** NGSPICE Simulation bench
.OPTION TUNING=FAST
.GLOBAL
** Default values that can be used or modified in the corners
.PARAM 
+ VDD=3.3 
+ VCM=1.65 
+ CL=6p 
+ IB=100u
+ VDD_MAX=3.63
+ VDD_MIN=2.97
+ T_MAX=75
+ T_MIN=0
.TEMP 27.0
**
** Process, Voltage and Temperature settings for nominal.
** Pyhton script replaces this include to simulate other corners
**
.lib "../../device_models/ptm130/ptm-130.lib" FNSP
.TEMP {T_MAX}
.PARAM vdd={VDD_MIN}
**
** Design variables for the circuit being simulated
**
.include 'design_var.inc'
*********** Unit Under Test ********************
.include "folded_cascode_ota.cir"
*********** Test-bench *************************
xi10 0 net15 vddnet vin vip vout folded_cascode_ota
c0 vout 0 cl
v2 vin 0 DC=vcm	
v1 vip 0 DC=vcm AC 1
v0 vddnet 0 DC=vdd
i1 vddnet net15 DC=100u

xi11 0 net16 vddd vinn vipp voutt folded_cascode_ota
c1 voutt 0 cl
v5 vipp 0 DC=vcm
v4 vinn 0 DC=vcm
v3 vddd 0 DC=vdd AC 1
i2 vddd net16 DC=100u
************************************************
** make params acessible in control
.csparam ib_sp = IB
.csparam cl_sp = CL
************************************************
.control
set units = degrees

let cl = $&cl_sp
print cl
AC DEC 21 1 1G
meas AC GDC FIND vdb(vout) at=1
meas AC GBW WHEN vdb(vout)=0
meas AC PM_Negative FIND vp(vout) WHEN vdb(vout)=0
meas AC GPS FIND vdb(voutt) at=1
let PM = PM_Negative + 180
let PSRR = GDC-GPS
print PM PSRR
************************************************
* Run noise
NOISE V(vout, 0) v1 dec 21 1 1G
print inoise_total onoise_total
let count = length(noise1.frequency)
echo "NOISE output $&count 3"
print noise1.all
OP
let idd = mag(i(v0)) - $&ib_sp
let outswing = 1.65 - @m.xi10.mnm6[vdsat] - @m.xi10.mnm8[vdsat]
print idd outswing 
let vov_mpm0 = @m.xi10.mpm0[vgs] - @m.xi10.mpm0[vth] 
let vov_mpm1 = @m.xi10.mpm1[vgs] - @m.xi10.mpm1[vth]
let vov_mpm3 = @m.xi10.mpm3[vgs] - @m.xi10.mpm3[vth]
let vov_mpm4 = @m.xi10.mpm4[vgs] - @m.xi10.mpm4[vth]
let vov_mpm5 = @m.xi10.mpm5[vgs] - @m.xi10.mpm5[vth]
let vov_mpm6 = @m.xi10.mpm6[vgs] - @m.xi10.mpm6[vth]
let vov_mnm1 = @m.xi10.mnm1[vgs] - @m.xi10.mnm1[vth] 
let vov_mnm2 = @m.xi10.mnm2[vgs] - @m.xi10.mnm2[vth] 
let vov_mnm3 = @m.xi10.mnm3[vgs] - @m.xi10.mnm3[vth] 
let vov_mnm4 = @m.xi10.mnm4[vgs] - @m.xi10.mnm4[vth] 
let vov_mnm5 = @m.xi10.mnm5[vgs] - @m.xi10.mnm5[vth] 
let vov_mnm6 = @m.xi10.mnm6[vgs] - @m.xi10.mnm6[vth] 
let vov_mnm7 = @m.xi10.mnm7[vgs] - @m.xi10.mnm7[vth] 
let vov_mnm8 = @m.xi10.mnm8[vgs] - @m.xi10.mnm8[vth] 
print vov_mpm0 vov_mpm1 vov_mpm3 vov_mpm4 vov_mpm5 vov_mpm6 vov_mnm1 vov_mnm2 vov_mnm3 vov_mnm4 vov_mnm5 vov_mnm6 vov_mnm7 vov_mnm8
let delta_mpm0 = @m.xi10.mpm0[vds] - @m.xi10.mpm0[vdsat]
let delta_mpm1 = @m.xi10.mpm1[vds] - @m.xi10.mpm1[vdsat]
let delta_mpm3 = @m.xi10.mpm3[vds] - @m.xi10.mpm3[vdsat]
let delta_mpm4 = @m.xi10.mpm4[vds] - @m.xi10.mpm4[vdsat]
let delta_mpm5 = @m.xi10.mpm5[vds] - @m.xi10.mpm5[vdsat]
let delta_mpm6 = @m.xi10.mpm6[vds] - @m.xi10.mpm6[vdsat]
let delta_mnm1 = @m.xi10.mnm1[vds] - @m.xi10.mnm1[vdsat]
let delta_mnm2 = @m.xi10.mnm2[vds] - @m.xi10.mnm2[vdsat]
let delta_mnm3 = @m.xi10.mnm3[vds] - @m.xi10.mnm3[vdsat]
let delta_mnm4 = @m.xi10.mnm4[vds] - @m.xi10.mnm4[vdsat]
let delta_mnm5 = @m.xi10.mnm5[vds] - @m.xi10.mnm5[vdsat]
let delta_mnm6 = @m.xi10.mnm6[vds] - @m.xi10.mnm6[vdsat]
let delta_mnm7 = @m.xi10.mnm7[vds] - @m.xi10.mnm7[vdsat]
let delta_mnm8 = @m.xi10.mnm8[vds] - @m.xi10.mnm8[vdsat]
print delta_mpm0 delta_mpm1 delta_mpm3 delta_mpm4 delta_mpm5 delta_mpm6 delta_mnm1 delta_mnm2 delta_mnm3 delta_mnm4 delta_mnm5 delta_mnm6 delta_mnm7 delta_mnm8

quit
.endc
.END
