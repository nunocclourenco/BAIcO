.include 'design_var.inc'

*********** Unit Under Test ********************
** Library name: amplificadores
** Cell name: nova_diff
** View name: schematic
.subckt AMP CMFB GND VBIASN VBIASP VDD VIN VIP VON VOP

mpm0 VOP net11 VDD VDD pch_lvt w='_wp0*_nfp0' l=_lp0 m=1 nf=_nfp0
mpm3 VON net41 VDD VDD pch_lvt w='_wp0*_nfp0' l=_lp0 m=1 nf=_nfp0
mpm1 net11 net11 VDD VDD pch_lvt w='_wp1*_nfp1' l=_lp1 m=1 nf=_nfp1
mpm2 net41 net41 VDD VDD pch_lvt w='_wp1*_nfp1' l=_lp1 m=1 nf=_nfp1
mpm5 vp VIN net26 VDD pch_lvt w='_wp5*_nfp5' l=_lp5 m=1 nf=_nfp5
mpm6 vn VIP net26 VDD pch_lvt w='_wp5*_nfp5' l=_lp5 m=1 nf=_nfp5
mpm4 net26 VBIASP VDD VDD pch_lvt w='_wp4*_nfp4' l=_lp4 m=1 nf=_nfp4
        
mnm0 net11 VIP vn GND nch_lvt l=_ln0 w='_wn0*_nfn0' m=1 nf=_nfn0
mnm1 net41 VIN vp GND nch_lvt l=_ln0 w='_wn0*_nfn0' m=1 nf=_nfn0
mnm5 VON CMFB GND GND nch_lvt l=_ln4 w='_wn4*_nfn4' m=1 nf=_nfn4
mnm4 VOP CMFB GND GND nch_lvt l=_ln4 w='_wn4*_nfn4' m=1 nf=_nfn4
mnm9 vn VBIASN GND GND nch_lvt l=_ln8 w='_wn8*_nfn8' m=1 nf=_nfn8
mnm8 vp VBIASN GND GND nch_lvt l=_ln8 w='_wn8*_nfn8' m=1 nf=_nfn8
mnm7 VDD VIN vn GND nch_lvt l=_ln6 w='_wn6*_nfn6' m=1 nf=_nfn6
mnm6 VDD VIP vp GND nch_lvt l=_ln6 w='_wn6*_nfn6' m=1 nf=_nfn6

.ends
************************************************