** NGSPICE Simulation bench

.GLOBAL
** Default values that can be modified in the corners
.PARAM vdd=3.3 vcm=1.65 c1=6p ib=100u
.TEMP 25.0
**
** Process, Voltage and Temperature settings for nominal.
** Pyhton script replaces this include to simulate other corners
**
.include 'nominal.corner'
**
** Design variables for the circuit being simulated
**
.include 'design_var.inc'

*********** Unit Under Test ********************
.include "ss_vc_ota.cir"

*********** Test-bench *************************
xmnmbias halfvdd halfvdd 0 0 nmos3v3 w='_w10/_nf10' l='_l10'  m='_nf10'
g2 cmfb 0 VCCS halfvdd 0 -1
g1 cmfb 0 VCCS outputn 0 -500m
g0 cmfb 0 VCCS outputp 0 -500m
e3 output 0 VCVS outputp outputn 1
i0 cmfb 0 DC 'vcm'
xinova cmfb 0 vddnet in_n in_p outputn outputp ss_vc_ota
cload2 outputp 0 'c1'
cload1 outputn 0 'c1'
r0 cmfb 0 1
cload3 output 0 'c1'
ibias vddnet halfvdd DC 'ib'
vin in_n 0 DC 'vcm'
vip in_p 0 DC 'vcm' AC 1 sin 'vcm' 100e-3 1e3
vdc vddnet 0 DC 'vdd'
************************************************

*********** OPTIONS ****************************
.OPTION KEEPOPINFO
************************************************


************************************************
** make params acessible in control
.csparam ib_sp = {ib}
.csparam cl_sp = {c1}
************************************************
.control
set units = degrees

***********************************************
** Run OP and save dc current, deltas and
** overdrives.

OP 
let idd = mag(i(vdc))  - $&ib_sp
print idd

let cl = $&cl_sp
print cl
** Overdrive and delta for  PMOS (in other simulator this is usualy defined inversly, but in ngspice it seems this is the way to go)
let vov_mpm0   = @m.xinova.xmpm0.xm1.msky130_fd_pr__pfet_g5v0d10v5[vgs] - @m.xinova.xmpm0.xm1.msky130_fd_pr__pfet_g5v0d10v5[vth] 
let delta_mpm0 = @m.xinova.xmpm0.xm1.msky130_fd_pr__pfet_g5v0d10v5[vds] - @m.xinova.xmpm0.xm1.msky130_fd_pr__pfet_g5v0d10v5[vdsat]
print vov_mpm0 delta_mpm0 

let   vov_mpm1 = @m.xinova.xmpm1.xm1.msky130_fd_pr__pfet_g5v0d10v5[vgs] - @m.xinova.xmpm1.xm1.msky130_fd_pr__pfet_g5v0d10v5[vth] 
let delta_mpm1 = @m.xinova.xmpm1.xm1.msky130_fd_pr__pfet_g5v0d10v5[vds] - @m.xinova.xmpm1.xm1.msky130_fd_pr__pfet_g5v0d10v5[vdsat]
print vov_mpm1 delta_mpm1 

let   vov_mpm2 = @m.xinova.xmpm2.xm1.msky130_fd_pr__pfet_g5v0d10v5[vgs] - @m.xinova.xmpm2.xm1.msky130_fd_pr__pfet_g5v0d10v5[vth] 
let delta_mpm2 = @m.xinova.xmpm2.xm1.msky130_fd_pr__pfet_g5v0d10v5[vds] - @m.xinova.xmpm2.xm1.msky130_fd_pr__pfet_g5v0d10v5[vdsat]
print vov_mpm2 delta_mpm2 

let   vov_mpm3 = @m.xinova.xmpm3.xm1.msky130_fd_pr__pfet_g5v0d10v5[vgs] - @m.xinova.xmpm3.xm1.msky130_fd_pr__pfet_g5v0d10v5[vth] 
let delta_mpm3 = @m.xinova.xmpm3.xm1.msky130_fd_pr__pfet_g5v0d10v5[vds] - @m.xinova.xmpm3.xm1.msky130_fd_pr__pfet_g5v0d10v5[vdsat]
print vov_mpm3 delta_mpm3 

** Overdrive and delta for NMOS
let   vov_mnm4 = @m.xinova.xmnm4.xm1.msky130_fd_pr__nfet_g5v0d10v5[vgs] - @m.xinova.xmnm4.xm1.msky130_fd_pr__nfet_g5v0d10v5[vth] 
let delta_mnm4 = @m.xinova.xmnm4.xm1.msky130_fd_pr__nfet_g5v0d10v5[vds] - @m.xinova.xmnm4.xm1.msky130_fd_pr__nfet_g5v0d10v5[vdsat]
print vov_mnm4 delta_mnm4

let   vov_mnm5 = @m.xinova.xmnm5.xm1.msky130_fd_pr__nfet_g5v0d10v5[vgs] - @m.xinova.xmnm5.xm1.msky130_fd_pr__nfet_g5v0d10v5[vth] 
let delta_mnm5 = @m.xinova.xmnm5.xm1.msky130_fd_pr__nfet_g5v0d10v5[vds] - @m.xinova.xmnm5.xm1.msky130_fd_pr__nfet_g5v0d10v5[vdsat]
print vov_mnm5 delta_mnm5

let   vov_mnm6 = @m.xinova.xmnm6.xm1.msky130_fd_pr__nfet_g5v0d10v5[vgs] - @m.xinova.xmnm6.xm1.msky130_fd_pr__nfet_g5v0d10v5[vth] 
let delta_mnm6 = @m.xinova.xmnm6.xm1.msky130_fd_pr__nfet_g5v0d10v5[vds] - @m.xinova.xmnm6.xm1.msky130_fd_pr__nfet_g5v0d10v5[vdsat]
print vov_mnm6 delta_mnm6

let   vov_mnm7 = @m.xinova.xmnm7.xm1.msky130_fd_pr__nfet_g5v0d10v5[vgs] - @m.xinova.xmnm7.xm1.msky130_fd_pr__nfet_g5v0d10v5[vth] 
let delta_mnm7 = @m.xinova.xmnm7.xm1.msky130_fd_pr__nfet_g5v0d10v5[vds] - @m.xinova.xmnm7.xm1.msky130_fd_pr__nfet_g5v0d10v5[vdsat]
print vov_mnm7 delta_mnm7

let   vov_mnm8 = @m.xinova.xmnm8.xm1.msky130_fd_pr__nfet_g5v0d10v5[vgs] - @m.xinova.xmnm8.xm1.msky130_fd_pr__nfet_g5v0d10v5[vth] 
let delta_mnm8 = @m.xinova.xmnm8.xm1.msky130_fd_pr__nfet_g5v0d10v5[vds] - @m.xinova.xmnm8.xm1.msky130_fd_pr__nfet_g5v0d10v5[vdsat]
print vov_mnm8 delta_mnm8

let   vov_mnm9 = @m.xinova.xmnm9.xm1.msky130_fd_pr__nfet_g5v0d10v5[vgs] - @m.xinova.xmnm9.xm1.msky130_fd_pr__nfet_g5v0d10v5[vth] 
let delta_mnm9 = @m.xinova.xmnm9.xm1.msky130_fd_pr__nfet_g5v0d10v5[vds] - @m.xinova.xmnm9.xm1.msky130_fd_pr__nfet_g5v0d10v5[vdsat]
print vov_mnm9 delta_mnm9

let   vov_mnm10 = @m.xinova.xmnm10.xm1.msky130_fd_pr__nfet_g5v0d10v5[vgs] - @m.xinova.xmnm10.xm1.msky130_fd_pr__nfet_g5v0d10v5[vth] 
let delta_mnm10 = @m.xinova.xmnm10.xm1.msky130_fd_pr__nfet_g5v0d10v5[vds] - @m.xinova.xmnm10.xm1.msky130_fd_pr__nfet_g5v0d10v5[vdsat]
print vov_mnm10 delta_mnm10

let   vov_mnm11 = @m.xinova.xmnm11.xm1.msky130_fd_pr__nfet_g5v0d10v5[vgs] - @m.xinova.xmnm11.xm1.msky130_fd_pr__nfet_g5v0d10v5[vth] 
let delta_mnm11 = @m.xinova.xmnm11.xm1.msky130_fd_pr__nfet_g5v0d10v5[vds] - @m.xinova.xmnm11.xm1.msky130_fd_pr__nfet_g5v0d10v5[vdsat]
print vov_mnm11 delta_mnm11
************************************************

************************************************
* Run AC
AC DEC 20 1 10G

let vdb_out = vdb(output)
let vp_out = vp(output)

let count = length(frequency)
echo "AC output $&count 3"
print frequency vdb_out vp_out


************************************************
* Run noise
NOISE V(output, 0) vip dec 20 0.01 10G
print inoise_total onoise_total
let count = length(noise2.frequency)
echo "NOISE output $&count 3"
print noise2.all

quit

.endc

.END
