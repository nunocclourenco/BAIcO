* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
.subckt  sky130_fd_pr__pfet_01v8 d g s b
+ 
.param  l = 1 w = 1 ad = 0 as = 0 pd = 0 ps = 0 nrd = 0 nrs = 0 sa = 0 sb = 0 sd = 0 mult = 1 nf = 1.0
msky130_fd_pr__pfet_01v8 d g s b sky130_fd_pr__pfet_01v8__model l = {l} w = {w} ad = {ad} as = {as} pd = {pd} ps = {ps} nrd = {nrd} nrs = {nrs} sa = {sa} sb = {sb} sd = {sd} nf = {nf}
.model sky130_fd_pr__pfet_01v8__model.0 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 7e-06 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.004443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.047954+0*(0.005856/sqrt(l*w*mult))}
+ k1 = 0.43448553
+ k2 = 0.022159346
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 160312.5
+ ua = -5.6628421e-10
+ ub = 1.06194446e-18
+ uc = -6.6549964e-11
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.011074
+ a0 = 1.198023
+ keta = 0.0051290095
+ a1 = 0.0
+ a2 = 0.9995
+ ags = 0.2608008
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.29454245+0*(0.0/sqrt(l*w*mult))}
+ nfactor = {1.5294758+0*(0.1/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.0015228006
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0029632464
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 9.3760948e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 4.6464006
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 1181082000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.4485
+ kt2 = -0.0075706
+ at = 90900.0
+ ute = -0.33954
+ ua1 = 1.6104e-9
+ ub1 = -5.609e-19
+ uc1 = -1.0858e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.1 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 7e-06 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.004443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.047954+0*(0.005856/sqrt(l*w*mult))}
+ k1 = 0.43448553
+ k2 = 0.022159346
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 160312.5
+ ua = -5.6628421e-10
+ ub = 1.06194446e-18
+ uc = -6.6549964e-11
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.011074
+ a0 = 1.198023
+ keta = 0.0051290095
+ a1 = 0.0
+ a2 = 0.9995
+ ags = 0.2608008
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.29454245+0*(0.0/sqrt(l*w*mult))}
+ nfactor = {1.5294758+0*(0.1/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.0015228006
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0029632464
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 9.3760948e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 4.6464006
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 1181082000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.4485
+ kt2 = -0.0075706
+ at = 90900.0
+ ute = -0.33954
+ ua1 = 1.6104e-9
+ ub1 = -5.609e-19
+ uc1 = -1.0858e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.2 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 7e-06 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.004443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.052801912332+0*(0.005856/sqrt(l*w*mult))} lvth0 = 3.8751001864043e-8
+ k1 = 0.438102126509735 lk1 = -2.89086783119324e-8
+ k2 = 0.021293418608066 lk2 = 6.92165032718695e-9
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 267009.4996875 lvsat = -0.852865182088082
+ ua = -5.79776770650915e-10 lua = 1.07850597768264e-16
+ ub = 1.0476535911495e-18 lub = 1.14231745035677e-25
+ uc = -7.3167975313894e-11 luc = 5.29000013197789e-17
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0108535677424 lu0 = 1.76198954109988e-9
+ a0 = 1.249119756379 la0 = -4.08433644441004e-7
+ keta = 0.0213163689759253 lketa = -1.29391035618573e-07 pketa = 5.04870979341448e-29
+ a1 = 0.0
+ a2 = 1.19866773275 la2 = -1.59201500656442e-6
+ ags = 0.22509732334312 lags = 2.85389956693552e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.306872589892495+0*(0.0/sqrt(l*w*mult))} lvoff = 9.85589757479963e-8
+ nfactor = {1.44269527408715+0*(0.1/sqrt(l*w*mult))} lnfactor = 6.9366607543917e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.429857606134414 lpclm = 3.44816939760565e-06 wpclm = 1.75362289861242e-22 ppclm = -1.40101696767252e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00576487163879899 lpdiblc2 = -2.2394337483051e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 1.01351357083584e-08 lpscbe2 = -6.06727053633572e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 3.2565334854499 lbeta0 = 1.11096776216837e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 8.4402431089145e-11 lagidl = 1.24676640282756e-16
+ bgidl = 1361862407.929 lbgidl = -1445.03890435438
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.43171925495647 lkt1 = -1.3413416702476e-7
+ kt2 = 0.0096543549776395 lkt2 = -1.37684887171055e-7
+ at = 87886.257761435 lat = 0.0240898603577266
+ ute = -0.47326335220418 lute = 1.06889595266106e-6
+ ua1 = 1.22719499268165e-09 lua1 = 3.06308714678805e-15
+ ub1 = -3.0164578823216e-19 lub1 = -2.07230654258392e-24
+ uc1 = -8.847741670786e-11 luc1 = -1.60686742927228e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.3 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 7e-06 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.004443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.053297910546+0*(0.005856/sqrt(l*w*mult))} lvth0 = 4.07316903799433e-8
+ k1 = 0.42438480066725 lk1 = 2.58692402332454e-8
+ k2 = 0.025136931386954 lk2 = -8.42679530623213e-9
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 53437.5
+ ua = -2.3668488550515e-10 lua = -1.26223126467596e-15
+ ub = 9.3695022895943e-19 lub = 5.56307687997067e-25
+ uc = -8.0533404316558e-11 luc = 8.2312648842419e-17
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0129883399648 lu0 = -6.76287749595451e-9
+ a0 = 1.168811571436 la0 = -8.77359177970925e-8
+ keta = -0.005560794812944 lketa = -2.20614361282578e-8
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.09661181618599 lags = 7.98476014873391e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.28931502304321+0*(0.0/sqrt(l*w*mult))} lvoff = 2.84456768612062e-8
+ nfactor = {1.6600217141216+0*(0.1/sqrt(l*w*mult))} lnfactor = -1.74191855955121e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.1592351855 leta0 = -3.16412877194199e-7
+ etab = -0.139268495071432 letab = 2.76612513571563e-7
+ dsub = 0.8590007 ldsub = -1.1940108573366e-6
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.46408247994329 lpclm = -1.21635517851718e-7
+ pdiblc1 = 0.39
+ pdiblc2 = -1.853824413469e-05 lpdiblc2 = 7.00772972043594e-10
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 800438663.92697 lpscbe1 = -1.75173332879876
+ pscbe2 = 8.2920612364473e-09 lpscbe2 = 1.29274878917682e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 3.9316215559846 lbeta0 = 8.41382277627077e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.3119513782171e-10 lagidl = -6.21824536352518e-17
+ bgidl = 918666228.2536 lbgidl = 324.793241398225
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.46634935213621 lkt1 = 4.15551598678871e-9
+ kt2 = -0.005808862085711 lkt2 = -7.5935034869729e-8
+ at = 106814.086142966 lat = -0.0514953559757196
+ ute = -0.17622069800093 lute = -1.17295765989642e-7
+ ua1 = 2.3392527360435e-09 lua1 = -1.37773529797308e-15
+ ub1 = -1.02790864263458e-18 lub1 = 8.27906511889728e-25
+ uc1 = -2.40574104777601e-10 luc1 = 4.46686741215816e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.4 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 7e-06 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.004443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.046167775834+0*(0.005856/sqrt(l*w*mult))} lvth0 = 2.65189219133937e-8
+ k1 = 0.3573341256955 lk1 = 1.59523898580084e-7
+ k2 = 0.052817427422536 lk2 = -6.36033799128071e-08 wk2 = -5.29395592033938e-23 pk2 = -5.04870979341448e-29
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 35743.666875 lvsat = 0.0352697899337212
+ ua = -7.6259585024292e-10 lua = -2.13912954047498e-16
+ ub = 1.15066129181608e-18 lub = 1.30309305384519e-25
+ uc = -4.286074864569e-11 luc = 7.21831273276241e-18
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0100904809916 lu0 = -9.86465086033959e-10
+ a0 = 1.282774495506 la0 = -3.1490254493694e-7
+ keta = -0.007016124315302 lketa = -1.91604725286866e-8
+ a1 = 0.0
+ a2 = 0.7006662 la2 = 1.980058382244e-7
+ ags = 0.3794348864849 lags = 2.34714041569902e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.2758638558486+0*(0.0/sqrt(l*w*mult))} lvoff = 1.6329541478367e-9
+ nfactor = {1.3656263388154+0*(0.1/sqrt(l*w*mult))} lnfactor = 4.12637632666988e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = -0.485738951 leta0 = 9.69238578108438e-07 weta0 = -1.32348898008484e-23 peta0 = 2.17725609840999e-28
+ etab = 7.38760593753566 letab = -1.47269923141726e-05 wetab = 1.79663629046518e-21 petab = -5.41158580981614e-28
+ dsub = 0.26
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.19003522874366 lpclm = 4.2463328176005e-7
+ pdiblc1 = 0.40797495771238 lpdiblc1 = -3.58301662564802e-8
+ pdiblc2 = 0.00023668464555664 lpdiblc2 = 1.92027487552058e-10
+ pdiblcb = -0.0490937606993659 lpdiblcb = 4.80270087649527e-8
+ drout = 0.40544946099372 ldrout = 3.080714623217e-7
+ pscbe1 = 799122672.14606 lpscbe1 = 0.871483095777194
+ pscbe2 = 8.9456362956796e-09 lpscbe2 = -1.00472122431867e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -4.4349697107106e-05 lalpha0 = 8.84041358658845e-11 walpha0 = -4.73671530539957e-27 palpha0 = -1.36295278593662e-32
+ alpha1 = 1.993338e-10 lalpha1 = -1.980058382244e-16
+ beta0 = -13.444963104552 lbeta0 = 4.30512292903355e-05 pbeta0 = 2.58493941422821e-26
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 807380539.7004 lbgidl = 546.623233247484
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.45647670127916 lkt1 = -1.55240141273016e-8
+ kt2 = -0.040468941952306 lkt2 = -6.84578058861025e-9
+ at = 71198.873273608 lat = 0.0194978012148608
+ ute = -0.16704404204188 lute = -1.35587943025743e-7
+ ua1 = 1.4237427767252e-09 lua1 = 4.47185493314543e-16
+ ub1 = -2.9305679836e-20 lub1 = -1.16264672076927e-24
+ uc1 = -2.1433991940186e-11 luc1 = 9.86642697270848e-18
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.5 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 7e-06 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.004443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.03759870481+0*(0.005856/sqrt(l*w*mult))} lvth0 = 1.8006938040556e-8
+ k1 = 0.55990344532888 lk1 = -4.16959042458991e-8
+ k2 = -0.032308223178728 lk2 = 2.09551636041513e-8
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 45098.15262 lvsat = 0.0259776237727545
+ ua = -6.248841862818e-10 lua = -3.50707182903309e-16
+ ub = 1.10184261276184e-18 lub = 1.788027543989e-25
+ uc = -5.7784011063288e-11 luc = 2.20421563761344e-17
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0109374520724 lu0 = -1.82779364549367e-9
+ a0 = 1.02077705376 la0 = -5.46505301478509e-8
+ keta = -0.0421967749919 lketa = 1.5785804653104e-8
+ a1 = 0.0
+ a2 = 0.9986676 la2 = -9.80102764488e-8
+ ags = 0.39549313889684 lags = 2.18762769235531e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.25992961562244+0*(0.0/sqrt(l*w*mult))} lvoff = -1.41951321699368e-8
+ nfactor = {1.9044637782592+0*(0.1/sqrt(l*w*mult))} lnfactor = -1.22610071755237e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.49
+ etab = -14.7771435475356 letab = 7.29009560982912e-6
+ dsub = 0.22117665755564 ldsub = 3.85647013369957e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.61200232157372 lpclm = 5.47733370242402e-9
+ pdiblc1 = 0.700518612109228 lpdiblc1 = -3.26424894827736e-7
+ pdiblc2 = 0.00043
+ pdiblcb = 0.220522721398732 lpdiblcb = -2.19793288329408e-07 wpdiblcb = -7.61006163548785e-23 ppdiblcb = 3.47098798297245e-29
+ drout = 0.43496363801256 ldrout = 2.7875390875016e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 8.7277890069796e-09 lpscbe2 = 2.06348777819499e-16
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 8.8699694214212e-05 lalpha0 = -4.37588804104509e-11
+ alpha1 = -9.86676e-11 lalpha1 = 9.80102764488e-17
+ beta0 = 50.1127373244192 lbeta0 = -2.00830497383779e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 1694552658.6996 lbgidl = -334.638545094944
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.43623405628508 lkt1 = -3.56318026204314e-8
+ kt2 = -0.03963756181126 lkt2 = -7.67162207515662e-9
+ at = 106443.99518944 lat = -0.015512517698768
+ ute = -0.23772148631908 lute = -6.53813518823178e-8
+ ua1 = 3.2739786116024e-09 lua1 = -1.39072407043071e-15
+ ub1 = -2.7909917868124e-18 lub1 = 1.58064103336246e-24 pub1 = 1.40129846432482e-45
+ uc1 = -4.6845503746344e-11 luc1 = 3.51086472872139e-17 puc1 = -1.17549435082229e-38
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.6 pmos
* DC IV MOS Parameters
+ lmin = 2.5e-07 lmax = 5e-07 wmin = 7e-06 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.006443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.990407688308+0*(0.007356/sqrt(l*w*mult))} lvth0 = -5.274183658508e-9
+ k1 = 0.13549433046384 lk1 = 1.6768123966339e-7
+ k2 = 0.11917144163576 lk2 = -5.37755112760986e-08 wk2 = -5.29395592033938e-23 pk2 = -6.31088724176809e-30
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 98492.4114752 lvsat = -0.000363793102352225
+ ua = -6.323516860368e-10 lua = -3.47023181509177e-16
+ ub = 1.1234768802288e-18 lub = 1.68129748155284e-25
+ uc = -2.5953323664251e-11 luc = 6.33886871606827e-18
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.01030450598072 lu0 = -1.51553728651644e-9
+ a0 = 1.15780283375864 la0 = -1.2225055440082e-7
+ keta = 0.059635137695792 lketa = -3.44517474884166e-08 wketa = -2.64697796016969e-23
+ a1 = 0.0
+ a2 = 0.8
+ ags = -0.33838723259592 lags = 5.80813843947026e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.22035128023192+0*(0.0/sqrt(l*w*mult))} lvoff = -3.37206289948251e-8
+ nfactor = {1.1039853562544+0*(0.1/sqrt(l*w*mult))} lnfactor = 2.72296351999767e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.965309351859001 leta0 = -2.34488165027416e-7
+ etab = 0.0047760499229952 letab = -2.38704054191061e-09 wetab = 2.68833699079734e-24 petab = -1.08468374467889e-30
+ dsub = 0.1852103104408 ldsub = 5.63082670899366e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.47758274175056 lpclm = 7.17916203732222e-8
+ pdiblc1 = -0.334384403489576 lpdiblc1 = 1.84132089081746e-07 wpdiblc1 = 2.11758236813575e-22 ppdiblc1 = 7.57306469012171e-29
+ pdiblc2 = -0.008973522524736 lpdiblc2 = 4.63911499530821e-09 wpdiblc2 = -4.96308367531817e-24 ppdiblc2 = -1.57772181044202e-30
+ pdiblcb = -0.3710028 lpdiblcb = 7.20287293464e-08 wpdiblcb = -4.2351647362715e-22
+ drout = 1.51703456660792 ldrout = -2.55072799021218e-7
+ pscbe1 = 800003445.66608 lpscbe1 = -0.00169987801257321
+ pscbe2 = 9.40358177202e-09 lpscbe2 = -1.27045473300003e-16
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -7.72393234514e-09 lalpha0 = 3.85984313528668e-15 walpha0 = -3.15544362088405e-30 palpha0 = -2.49204802374325e-36
+ alpha1 = 1.973352e-10 lalpha1 = -4.80191528976e-17
+ beta0 = 3.3812716986096 lbeta0 = 2.97135805052774e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 484651822.7312 lbgidl = 262.251513520035
+ cgidl = 527.777841138384 lcgidl = -0.000112371464591528
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.45936412512 lkt1 = -2.42208607215494e-8
+ kt2 = 0.00980465974399998 lkt2 = -3.20633487727855e-08 pkt2 = -2.52435489670724e-29
+ at = 63319.776 lat = 0.005762298347712
+ ute = -0.377306802 lute = 3.481388585076e-9
+ ua1 = 7.667833132e-10 lua1 = -1.53829356307462e-16 wua1 = 7.88860905221012e-31 pua1 = 1.88079096131566e-37
+ ub1 = 4.3271957856e-19 lub1 = -9.73828420763331e-27
+ uc1 = 1.101914492e-11 luc1 = 6.56181724345704e-18
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.24e-6
+ sbref = 1.24e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.7 pmos
* DC IV MOS Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 7e-06 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.006443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.790897759485714+0*(0.007356/sqrt(l*w*mult))} lvth0 = -5.38225307182653e-8
+ k1 = 0.335246697368572 lk1 = 1.19073898205527e-7
+ k2 = 0.0606923753943428 lk2 = -3.95453322550446e-8
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 158397.929237143 lvsat = -0.0149410819835079
+ ua = -1.56074952462286e-09 lua = -1.21108708263323e-16
+ ub = 1.39430136593714e-18 lub = 1.02227859451988e-25
+ uc = -4.91771559457713e-14 luc = 3.54055130302881e-20
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.00571223023114286 lu0 = -3.9806209016584e-10
+ a0 = 0.962178920290572 la0 = -7.46478225453271e-8
+ keta = -0.226972829022943 lketa = 3.52908619169869e-8
+ a1 = 0.0
+ a2 = 0.870068692128286 la2 = -1.70503754051129e-8
+ ags = 4.02569816488 lags = -4.81133968503969e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.149163822694+0*(0.0/sqrt(l*w*mult))} lvoff = -5.10432425371874e-8
+ nfactor = {0.604458806285715+0*(0.1/sqrt(l*w*mult))} lnfactor = 3.93850143616047e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = -0.417167463843577 leta0 = 1.01920978352018e-07 weta0 = -1.12496563307212e-22
+ etab = 0.124203059314531 letab = -3.14481701532282e-08 petab = 3.15544362088405e-30
+ dsub = 0.747409855918 ldsub = -8.04962459073943e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.10997007392457 lpclm = -8.20922482633373e-8
+ pdiblc1 = 1.00596961163057 lpdiblc1 = -1.4202697624956e-07 wpdiblc1 = 1.6940658945086e-21
+ pdiblc2 = 0.0247436758567886 lpdiblc2 = -3.56556062445522e-9
+ pdiblcb = -0.075
+ drout = -0.722076222894571 ldrout = 2.89787942274739e-7
+ pscbe1 = 799987694.049715 lpscbe1 = 0.00213308881063767
+ pscbe2 = 8.09092591147142e-09 lpscbe2 = 1.92373578494165e-16
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.80426155183571e-08 lalpha0 = -4.84351708872099e-15
+ alpha1 = -2.47625714285714e-10 lalpha1 = 6.02567460628571e-17
+ beta0 = 32.89328272192 lbeta0 = -4.21003568786257e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 6.77947653402857e-11 lagidl = 7.83675739162556e-18
+ bgidl = 2954967410.85428 lbgidl = -338.87014106266
+ cgidl = -513.492289779943 lcgidl = 0.000141009126525876 wcgidl = -2.16840434497101e-19
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.5589
+ kt2 = -0.12196
+ at = 208336.6 lat = -0.0295258055708
+ ute = -0.5190042 lute = 3.79617500196e-8
+ ua1 = 1.3462e-10
+ ub1 = 3.927e-19
+ uc1 = 3.7985e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.8 pmos
* DC IV MOS Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 7e-06 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.006443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.711113737733333+0*(0.007356/sqrt(l*w*mult))} lvth0 = -6.76521334807794e-8
+ k1 = -0.249508425106668 lk1 = 2.20434181625139e-7
+ k2 = 0.343856885470667 lk2 = -8.86285021026544e-8
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 197157.557086667 lvsat = -0.0216595983556886
+ ua = -9.60007983346665e-10 lua = -2.25240045545056e-16
+ ub = 6.24599095426667e-19 lub = 2.35646511617732e-25
+ uc = 2.69835080537333e-13 luc = -1.98914300172203e-20
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.00603241996793333 lu0 = -4.53563138761628e-10
+ a0 = -0.791160669612 la0 = 2.29272555289205e-7
+ keta = -0.0915648642361733 lketa = 1.18195161167778e-8
+ a1 = 0.0
+ a2 = -0.316691314966 la2 = 1.88660230704597e-7
+ ags = 1.25
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.390263853465334+0*(0.0/sqrt(l*w*mult))} lvoff = -9.25144540334603e-9
+ nfactor = {-0.669046547333334+0*(0.1/sqrt(l*w*mult))} lnfactor = 6.14597014601666e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = -0.617243906024667 leta0 = 1.36601828686804e-7
+ etab = -0.246957641957333 letab = 3.28880834838343e-8
+ dsub = 0.393013456590667 ldsub = -1.9065882840793e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.11806085162867 lpclm = -2.5683268748901e-07 wpclm = 3.3881317890172e-21
+ pdiblc1 = 0.985023109708667 lpdiblc1 = -1.38396151499421e-7
+ pdiblc2 = 0.0220607773736267 lpdiblc2 = -3.1005123671809e-9
+ pdiblcb = -0.418610236790253 lpdiblcb = 5.95607112247489e-8
+ drout = 0.709556465021333 ldrout = 4.16315954167721e-8
+ pscbe1 = 867303832.327334 lpscbe1 = -11.6663116879553
+ pscbe2 = 1.013312288888e-08 lpscbe2 = -1.61616761175883e-16
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 14.4732975792 lbeta0 = -1.01715230319377e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.75145547539333e-10 lagidl = -1.0771212493193e-17
+ bgidl = 780957079.713333 lbgidl = 37.9684617166503
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = 0.0674870599999995 lkt1 = -1.0857668020628e-7
+ kt2 = -0.12196
+ at = 38000.0
+ ute = -0.3
+ ua1 = 1.3462e-10
+ ub1 = 3.927e-19
+ uc1 = 3.7985e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.9 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.004443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.062648749802+0*(0.005856/sqrt(l*w*mult))} wvth0 = 1.03594197797603e-7
+ k1 = 0.444388049205489 wk1 = -6.98102075292465e-8
+ k2 = 0.0180906853887137 wk2 = 2.86830084088628e-8
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 160312.5
+ ua = -5.9463144281392e-10 wua = 1.99840683421517e-16
+ ub = 1.01974565808793e-18 wub = 2.97490674628997e-25
+ uc = -7.49378332315679e-11 wuc = 5.91323156898652e-17
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.01117524733111 wu0 = -7.13767582763556e-10
+ a0 = 1.2066858327441 wa0 = -6.10707375676198e-8
+ keta = 0.0303539152578079 wketa = -1.77829082611841e-7
+ a1 = 0.0
+ a2 = 1.22604688730313 wa2 = -1.59709715169954e-6
+ ags = 0.343036381949931 wags = -5.79739652413986e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.306629209945388+0*(0.0/sqrt(l*w*mult))} wvoff = 8.52085416482716e-8
+ nfactor = {1.06134045929744+0*(0.1/sqrt(l*w*mult))} wnfactor = 3.30023346666222e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.56849442030249 wpclm = 4.018474456923e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0100191156662281 wpdiblc2 = -4.9742059323811e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 1.01311090249299e-08 wpscbe2 = -5.32265564308848e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 0.342093011489364 wbeta0 = 3.03442588485037e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 268797089.07066 wbgidl = 6431.37343500181
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.479925454664196 wkt1 = 2.21541353900369e-7
+ kt2 = 0.100910653452993 wkt2 = -7.64764870376458e-7
+ at = 93172.3839899999 wat = -0.0160197213089073
+ ute = -0.780957886934979 wute = 3.11188230536035e-6
+ ua1 = 7.2932880804441e-10 wua1 = 6.21132476313363e-15
+ ub1 = -7.73186088509244e-20 wub1 = -3.40912414031835e-24
+ uc1 = -6.65340992675926e-10 wuc1 = 3.92502146538137e-15
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.10 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.004443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.062648749802+0*(0.005856/sqrt(l*w*mult))} wvth0 = 1.03594197797603e-7
+ k1 = 0.444388049205489 wk1 = -6.98102075292448e-8
+ k2 = 0.0180906853887137 wk2 = 2.86830084088628e-8
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 160312.5
+ ua = -5.94631442813919e-10 wua = 1.99840683421519e-16
+ ub = 1.01974565808792e-18 wub = 2.97490674628997e-25
+ uc = -7.49378332315677e-11 wuc = 5.91323156898654e-17
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.01117524733111 wu0 = -7.13767582763556e-10
+ a0 = 1.2066858327441 wa0 = -6.10707375676232e-8
+ keta = 0.0303539152578079 wketa = -1.77829082611841e-7
+ a1 = 0.0
+ a2 = 1.22604688730313 wa2 = -1.59709715169953e-6
+ ags = 0.343036381949931 wags = -5.79739652413987e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.306629209945388+0*(0.0/sqrt(l*w*mult))} wvoff = 8.52085416482716e-8
+ nfactor = {1.06134045929744+0*(0.1/sqrt(l*w*mult))} wnfactor = 3.30023346666222e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.56849442030249 wpclm = 4.018474456923e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0100191156662281 wpdiblc2 = -4.9742059323811e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 1.01311090249299e-08 wpscbe2 = -5.32265564308848e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 0.342093011489364 wbeta0 = 3.03442588485036e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 268797089.070658 wbgidl = 6431.37343500181
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.479925454664195 wkt1 = 2.21541353900371e-7
+ kt2 = 0.100910653452993 wkt2 = -7.64764870376458e-7
+ at = 93172.3839899999 wat = -0.0160197213089077
+ ute = -0.780957886934979 wute = 3.11188230536035e-6
+ ua1 = 7.29328808044408e-10 wua1 = 6.21132476313363e-15
+ ub1 = -7.73186088509237e-20 wub1 = -3.40912414031835e-24
+ uc1 = -6.65340992675926e-10 wuc1 = 3.92502146538137e-15
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.11 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.004443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.06298214945842+0*(0.005856/sqrt(l*w*mult))} lvth0 = 2.66497614281229e-09 wvth0 = 7.17680472761011e-08 pvth0 = 2.5439717835725e-13
+ k1 = 0.417739211580813 lk1 = 2.13013166441158e-07 wk1 = 1.43553300689437e-07 pk1 = -1.70548663805771e-12
+ k2 = 0.0275206297122963 lk2 = -7.53767322995775e-08 wk2 = -4.39002329098013e-08 pk2 = 5.80182380995648e-13
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 275393.831959135 lvsat = -0.919883983839571 wvsat = -0.0591073810341687 pvsat = 4.72465274900901e-7
+ ua = -2.51490382696535e-10 lua = -2.74284247519658e-15 wua = -2.31433440284757e-15 pua = 2.0096651255728e-20
+ ub = 7.43366684165797e-19 lub = 2.20919055465276e-24 wub = 2.14514424907052e-24 pub = -1.47689195274193e-29
+ uc = -9.31427811835541e-11 luc = 1.45518302252635e-16 wuc = 1.40817231876151e-16 puc = -6.52935144578655e-22
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.01215566032122 lu0 = -7.83677240953952e-09 wu0 = -9.17941700121389e-09 pu0 = 6.76687971911769e-14
+ a0 = 1.35606158915781 la0 = -1.19401091002048e-06 wa0 = -7.53912351486146e-07 pa0 = 5.53811720051629e-12
+ keta = 0.0733454834213588 lketa = -3.43646135481302e-07 wketa = -3.66791843734603e-07 pketa = 1.51044321906749e-12
+ a1 = 0.0
+ a2 = 1.65138419351546 la2 = -3.39986485256465e-06 wa2 = -3.19153433809292e-06 pa2 = 1.27448753506113e-11
+ ags = 0.418601350570406 lags = -6.0401633514285e-07 wags = -1.36415350661415e-06 pags = 6.27008506850459e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.347588216412412+0*(0.0/sqrt(l*w*mult))} lvoff = 3.27399182835104e-07 wvoff = 2.87034670476895e-07 pvoff = -1.61326446495874e-12
+ nfactor = {0.583466011452519+0*(0.1/sqrt(l*w*mult))} lnfactor = 3.81981198318783e-06 wnfactor = 6.05734479227026e-06 pnfactor = -2.20385227292131e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -1.55231284286998 lpclm = 7.86399318220881e-06 wpclm = 7.91302005002574e-06 ppclm = -3.11304192820806e-11
+ pdiblc1 = 0.39
+ pdiblc2 = 0.019740218572311 lpdiblc2 = -7.77040612611031e-08 wpdiblc2 = -9.85225930368203e-08 ppdiblc2 = 3.89919293788478e-13
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 1.37853598461252e-08 lpscbe2 = -2.92096619505918e-14 wpscbe2 = -2.57331391434733e-14 ppscbe2 = 1.63147893361998e-19
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = -3.75323786342985 lbeta0 = 3.27353639050649e-05 wbeta0 = 4.94170808905484e-05 pbeta0 = -1.52455513195914e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 4.50205801158688e-11 lagidl = 4.39469086177782e-16 wagidl = 2.77631896720417e-16 pagidl = -2.21920559006739e-21
+ bgidl = 765453235.265036 lbgidl = -3969.94044630906 wbgidl = 4204.53091299624 pbgidl = 0.017799904951163
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.488364753628569 lkt1 = 6.74581691052819e-08 wkt1 = 3.99336162428739e-07 pkt1 = -1.42117399921254e-12
+ kt2 = 0.159378129288713 lkt2 = -4.67350296361748e-07 wkt2 = -1.05551401010405e-06 pkt2 = 2.3240561470519e-12
+ at = 93442.9686279172 lat = -0.00216287446848007 wat = -0.0391733790886386 pat = 1.85075012569723e-7
+ ute = -1.35535786977856 lute = 4.59137321006297e-06 wute = 6.21853894493278e-06 pute = -2.48325565700466e-11
+ ua1 = -6.18676573154753e-11 lua1 = 6.32430077202686e-15 wua1 = 9.08755936212857e-15 pua1 = -2.2990715317061e-20
+ ub1 = 4.06081585772902e-19 lub1 = -3.86398114489403e-24 wub1 = -4.98929553461867e-24 pub1 = 1.26308440525738e-29
+ uc1 = -1.20516963553766e-09 luc1 = 4.31503280447514e-15 wuc1 = 7.87239225949609e-15 puc1 = -3.15526689686874e-20
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.12 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.004443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.07636237298153+0*(0.005856/sqrt(l*w*mult))} lvth0 = 5.60967311861451e-08 wvth0 = 1.6259851415204e-07 pvth0 = -1.08319576576196e-13
+ k1 = 0.516176246160522 lk1 = -1.80079184353312e-07 wk1 = -6.47106026892919e-07 pk1 = 1.45188329983136e-12
+ k2 = -0.00637185451196262 lk2 = 5.99674128675563e-08 wk2 = 2.22128817622357e-07 pk2 = -4.82161535598342e-13
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 36668.8354567295 lvsat = 0.0334256162433536 wvsat = 0.118214762068338 pvsat = -2.35641977391776e-7
+ ua = -1.2930637317316e-09 lua = 1.41651195929239e-15 wua = 7.44719853142989e-15 pua = -1.88844491489737e-20
+ ub = 1.51150319542223e-18 lub = -8.58238164935004e-25 wub = -4.05045029380802e-24 pub = 9.97218359325022e-30
+ uc = -6.19625728364736e-11 luc = 2.10051914123208e-17 wuc = -1.30919574374239e-16 puc = 4.32201769819667e-22
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.00925930203023656 lu0 = 3.72936521545947e-09 wu0 = 2.62887560926926e-08 pu0 = -7.39676062152977e-14
+ a0 = 1.13431230231456 la0 = -3.08491056396393e-07 wa0 = 2.43210953394609e-07 pa0 = 1.55626681645033e-12
+ keta = -0.00909786835714493 lketa = -1.44219659768352e-08 wketa = 2.4935456629057e-08 pketa = -5.38562951121243e-14
+ a1 = 0.0
+ a2 = 0.8
+ ags = -0.112013842866754 lags = 1.51490948018711e-06 wags = 1.47075711262695e-06 pags = -5.0506712339144e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.293835593771702+0*(0.0/sqrt(l*w*mult))} lvoff = 1.12746792244301e-07 wvoff = 3.18688582327384e-08 pvoff = -5.94301130623276e-13
+ nfactor = {1.33820912601027+0*(0.1/sqrt(l*w*mult))} lnfactor = 8.05867623585996e-07 wnfactor = 2.26869578289966e-06 pnfactor = -6.90916667143107e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.15923519030644 leta0 = -3.16412896387939e-07 weta0 = -3.38841630738418e-14 peta0 = 1.35310916267557e-19
+ etab = -0.139268495046268 letab = 2.76612513471073e-07 wetab = -1.77403851022362e-16 petab = 7.08434150418352e-22
+ dsub = 0.8590007 ldsub = -1.1940108573366e-6
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.02474689264385 lpclm = -2.42707738788853e-06 wpclm = -3.95253957025334e-06 ppclm = 1.62527708408454e-11
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00047479002903789 lpdiblc2 = -7.70693372965986e-10 wpdiblc2 = -3.47783714583786e-09 ppdiblc2 = 1.03734583882938e-14
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 772483502.723579 lpscbe1 = 109.882674200826 wpscbe1 = 197.076679643345 ppscbe1 = -0.000786993793733592
+ pscbe2 = 5.30349045775227e-09 lpscbe2 = 4.66130938903466e-15 wpscbe2 = 2.10686535362533e-14 ppscbe2 = -2.37474838140749e-20
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 0.949781421168005 lbeta0 = 1.39546182811475e-05 wbeta0 = 2.10212042320702e-05 pbeta0 = -3.90611798923001e-11
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 2.09958839768263e-10 lagidl = -2.19185133745989e-16 wagidl = -5.55263793440834e-16 pagidl = 1.10682841948977e-21
+ bgidl = -871227871.615888 lbgidl = 2565.8804116806 wbgidl = 12618.291969381 pbgidl = -0.0157990867982182
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.481238919034349 lkt1 = 3.90023030384709e-08 wkt1 = 1.04967608101537e-07 pkt1 = -2.45660865212659e-13
+ kt2 = 0.126050459846816 lkt2 = -3.34261647527979e-07 wkt2 = -9.29574226291119e-07 pkt2 = 1.82113602263992e-12
+ at = 101167.433209994 lat = -0.0330092724137401 wat = 0.0398074474703289 pat = -1.30322123399613e-7
+ ute = -0.326436011397087 lute = 4.82540453957603e-07 wute = 1.05897923393512e-06 pute = -4.22869071285058e-12
+ ua1 = 1.02204857932899e-09 lua1 = 1.99585687541753e-15 wua1 = 9.28594972960573e-15 pua1 = -2.37829551103415e-20
+ ub1 = -3.50091720583559e-19 lub1 = -8.44325546035128e-25 wub1 = -4.7784345592572e-24 pub1 = 1.17888049069457e-29
+ uc1 = 9.61647670837893e-11 luc1 = -8.81635316220402e-16 wuc1 = -2.37392223534164e-15 puc1 = 9.36432806349893e-21
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.13 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.004443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.06309909752088+0*(0.005856/sqrt(l*w*mult))} lvth0 = 2.96585402059754e-08 wvth0 = 1.19361452997798e-07 pvth0 = -2.21334995691011e-14
+ k1 = 0.327480830921503 lk1 = 1.96054557268403e-07 wk1 = 2.10458031977282e-07 pk1 = -2.57531726148844e-13
+ k2 = 0.0589027282408705 lk2 = -7.01468933678106e-08 wk2 = -4.28998019787076e-08 pk2 = 4.61300829400061e-14
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -72820.2721227911 lvsat = 0.2516744149677 wvsat = 0.765347782150954 pvsat = -1.52559681737722e-6
+ ua = -5.76104297463658e-10 lua = -1.26305254923907e-17 wua = -1.31471736957148e-15 pua = -1.41898923070343e-21
+ ub = 1.06757465867557e-18 lub = 2.66614566465191e-26 wub = 5.85739343906578e-25 pub = 7.30690613187482e-31
+ uc = -5.36881133222912e-11 luc = 4.51139683323947e-18 wuc = 7.63301296754247e-17 puc = 1.90830592487178e-23
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0111350245963138 lu0 = -9.58385295977659e-12 wu0 = -7.36376312989099e-09 pu0 = -6.88676085319117e-15
+ a0 = 0.213430063358942 la0 = 1.52713850403891e-06 wa0 = 7.53860256964215e-06 pa0 = -1.29859145170973e-11
+ keta = -0.0713723724377544 lketa = 1.09712169438199e-07 wketa = 4.53694958222524e-07 pketa = -9.08518902499442e-13
+ a1 = 0.0
+ a2 = 0.44986115912682 la2 = 6.97945056788462e-07 wa2 = 1.76811088061638e-06 pa2 = -3.52444260654609e-12
+ ags = 2.16149251083439 lags = -3.01695712788683e-06 wags = -1.25630468372084e-05 pags = 2.29234434638425e-11
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.22592411111109+0*(0.0/sqrt(l*w*mult))} lvoff = -2.26237467794384e-08 wvoff = -3.52062325933252e-07 pvoff = 1.71003488159794e-13
+ nfactor = {1.65671111183595+0*(0.1/sqrt(l*w*mult))} lnfactor = 1.70985512164207e-07 wnfactor = -2.05207260814041e-06 pnfactor = 1.70358515162794e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = -0.48573896061288 leta0 = 9.69238587657277e-07 weta0 = 6.77683260219522e-14 peta0 = -6.73168551339275e-20
+ etab = 26.0397399007306 letab = -5.190699972415e-05 wetab = -0.000131492735920389 petab = 2.6210946723443e-10
+ dsub = 0.26
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -1.49136427670448 lpclm = 2.58838261819793e-06 wpclm = 1.18534330486169e-05 ppclm = -1.52538750073081e-11
+ pdiblc1 = 0.431440277336474 lpdiblc1 = -8.26044795453339e-08 wpdiblc1 = -1.65424453990468e-07 ppdiblc1 = 3.29746850268454e-13
+ pdiblc2 = -0.000251411706063657 lpdiblc2 = 6.7687214127786e-10 wpdiblc2 = 3.44095344768364e-09 ppdiblc2 = -3.41802981581517e-15
+ pdiblcb = -0.0491388386668577 lpdiblcb = 4.81168643905167e-08 wpdiblcb = 3.17788049716879e-10 ppdiblcb = -6.33458995446526e-16
+ drout = 0.646986001581431 ldrout = -1.73392502420327e-07 wdrout = -1.7027703430232e-06 pdrout = 3.39419683002118e-12
+ pscbe1 = 855032994.55284 lpscbe1 = -54.6663647431296 wpscbe1 = -394.153359286687 ppscbe1 = 0.00039152750960712
+ pscbe2 = 2.02894901206716e-09 lpscbe2 = 1.11885772852937e-14 wpscbe2 = 4.8760862227486e-14 ppscbe2 = -7.89474157022394e-20
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -0.000156327218113701 lalpha0 = 3.11613183634129e-10 walpha0 = 7.89412655291583e-10 palpha0 = -1.57356624347361e-15
+ alpha1 = 4.5013884087318e-10 lalpha1 = -6.97945056788463e-16 walpha1 = -1.76811088061638e-15 palpha1 = 3.5244426065461e-21
+ beta0 = -66.4278004856646 lbeta0 = 0.000148260912644149 wbeta0 = 0.000373515344561367 pbeta0 = -7.4170114458802e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = -956458108.46995 lbgidl = 2735.7730815508 wbgidl = 12434.6077519975 pbgidl = -0.0154329420677075
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.456094110366761 lkt1 = -1.11197995813612e-08 wkt1 = -2.69716730047349e-09 pkt1 = -3.10485771423662e-14
+ kt2 = -0.036836989935945 lkt2 = -9.57190415291038e-09 wkt2 = -2.56043253981149e-08 pkt2 = 1.92184683336611e-14
+ at = -85625.6790834141 lat = 0.339332536458977 wat = 1.10557266474741 pat = -2.25475243007627e-6
+ ute = 0.292903058864427 lute = -7.52011649679342e-07 wute = -3.24250848702685e-06 pute = 4.3456282178763e-12
+ ua1 = 2.24902479407497e-09 lua1 = -4.49921438531804e-16 wua1 = -5.81802546461183e-15 pua1 = 6.32437259534972e-21
+ ub1 = -4.44619375295072e-19 lub1 = -6.55899979847783e-25 wub1 = 2.92785448511578e-24 pub1 = -3.57243388418665e-30
+ uc1 = -6.77736364354485e-10 luc1 = 6.61011217318505e-16 wuc1 = 4.6267625307692e-15 puc1 = -4.59040290681092e-21
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.14 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.004443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.02004338370715+0*(0.005856/sqrt(l*w*mult))} lvth0 = -1.31103364423258e-08 wvth0 = -1.2376048801328e-07 pvth0 = 2.19368763070956e-13
+ k1 = 0.5888156193584 lk1 = -6.35392188079261e-08 wk1 = -2.03823373349649e-07 pk1 = 1.53989736455796e-13
+ k2 = -0.0346694007439822 lk2 = 2.2801858093745e-08 wk2 = 1.66456931234654e-08 pk2 = -1.30187200737962e-14
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 184285.666797988 lvsat = -0.00371868418798851 wvsat = -0.98123609241366 pvsat = 2.09351315415046e-7
+ ua = 1.28371693700096e-10 lua = -7.12413297603014e-16 wua = -5.31025976450652e-15 pua = 2.54993486079655e-21
+ ub = 6.4775416056259e-19 lub = 4.4368511060107e-25 wub = 3.20120652400173e-24 pub = -1.86735232455388e-30
+ uc = -8.17040323518775e-11 luc = 3.23406738102506e-17 wuc = 1.68629983503067e-16 puc = -7.2601892952725e-23
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0145941945291977 lu0 = -3.44570879575081e-09 wu0 = -2.57790916122185e-08 pu0 = 1.14058847107871e-14
+ a0 = 2.56128558840139 la0 = -8.05075607495703e-07 wa0 = -1.08601880261215e-05 pa0 = 5.29030333571741e-12
+ keta = 0.0783135022673772 lketa = -3.89764979696472e-08 wketa = -8.49566387128427e-07 pketa = 3.8606011576878e-13
+ a1 = 0.0
+ a2 = 1.50658462837287 la2 = -3.51738520705474e-07 wa2 = -3.58068410901885e-06 pa2 = 1.78871871086818e-12
+ ags = -2.44917447063237 lags = 1.5629935901494e-06 wags = 2.00541732918712e-05 pags = -9.47648074473716e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.225907583557786+0*(0.0/sqrt(l*w*mult))} lvoff = -2.26401642261826e-08 wvoff = -2.39846555175946e-07 pvoff = 5.95352988672683e-14
+ nfactor = {2.5391686126243+0*(0.1/sqrt(l*w*mult))} lnfactor = -7.05593056753885e-07 wnfactor = -4.47450545536764e-06 pnfactor = 4.10987975122694e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.49
+ etab = -52.0813336230975 letab = 2.56936312078623e-05 wetab = 0.00026298492301251 petab = -1.29740181534657e-10
+ dsub = 0.202823170331954 ldsub = 5.67959176287979e-08 wdsub = 1.29387353397984e-07 pdsub = -1.28525374849646e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.60098323812158 lpclm = -4.83363677484353e-07 wpclm = -6.97206050238212e-06 ppclm = 3.4462031056541e-12
+ pdiblc1 = 0.605375734770895 lpdiblc1 = -2.55381178962326e-07 wpdiblc1 = 6.70732757401469e-07 ppdiblc1 = -5.0083988178119e-13
+ pdiblc2 = 0.00043
+ pdiblcb = 0.220612877333715 lpdiblcb = -2.19837765678061e-07 wpdiblcb = -6.35576099433757e-10 ppdiblcb = 3.13553841742194e-16
+ drout = -0.048109443162863 ldrout = 5.17072216471081e-07 wdrout = 3.40554068604641e-06 pdrout = -1.68008263097276e-12
+ pscbe1 = 800000000.0
+ pscbe2 = -2.90988437955433e-09 lpscbe2 = 1.60945081688602e-14 wpscbe2 = 8.20425971828652e-14 ppscbe2 = -1.12007427739346e-19
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.000312654736227403 lalpha0 = -1.54244412927155e-10 walpha0 = -1.57882531058317e-09 palpha0 = 7.78894521072479e-16
+ alpha1 = -6.0027768174636e-10 lalpha1 = 3.45473590957386e-16 walpha1 = 3.53622176123277e-15 palpha1 = -1.74455257124305e-21
+ beta0 = 155.296247045962 lbeta0 = -7.19860092828218e-05 wbeta0 = -0.000741516627228073 pbeta0 = 3.65902484205359e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 3074764530.63407 lbgidl = -1268.59355233152 wbgidl = -9730.13787851747 pbgidl = 0.00658414202741697
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.426665543009719 lkt1 = -4.03523138226714e-08 wkt1 = -6.74555518285744e-08 pkt1 = 3.32783870280045e-14
+ kt2 = -0.0378742970358044 lkt2 = -8.54150759295034e-09 wkt2 = -1.24305620973031e-08 pkt2 = 6.13246864395923e-15
+ at = 424290.024863283 lat = -0.167186109068027 wat = -2.24073256849414 pat = 1.06925971770142e-6
+ ute = -0.425714525253207 lute = -3.81814959071009e-08 wute = 1.32530245988015e-06 pute = -1.91751972502409e-13
+ ua1 = 3.09442042783544e-09 lua1 = -1.28968504658016e-15 wua1 = 1.26583890545727e-15 pua1 = -7.12299070285965e-22
+ ub1 = -2.5174169121692e-18 lub1 = 1.40308857983569e-24 wub1 = -1.92863233863185e-24 pub1 = 1.25169902434118e-30
+ uc1 = -4.84160950733e-11 luc1 = 3.58834796712717e-17 wuc1 = 1.10722639565959e-17 puc1 = -5.46236855581912e-24
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.15 pmos
* DC IV MOS Parameters
+ lmin = 2.5e-07 lmax = 5e-07 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.006443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.08819162925908+0*(0.007356/sqrt(l*w*mult))} lvth0 = 2.05097827217694e-08 wvth0 = 6.89351575005131e-07 pvth0 = -1.81770315874422e-13
+ k1 = 0.102010233858814 lk1 = 1.76620376463669e-07 wk1 = 2.36054248865334e-07 pk1 = -6.30186099324991e-14
+ k2 = 0.126991335773725 lk2 = -5.69515263384275e-08 wk2 = -5.51282377039432e-08 pk2 = 2.23900874127359e-14
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 214586.750038586 lvsat = -0.0186673599917385 wvsat = -0.818435157751386 pvsat = 1.29035427910629e-7
+ ua = -5.57954408339692e-10 lua = -3.7382255107491e-16 wua = -5.24481628146432e-16 pua = 1.88928646560936e-22
+ ub = 1.34258818152846e-18 lub = 1.00897084365813e-25 wub = -1.54467818726909e-24 pub = 4.73972947135051e-31
+ uc = -3.19062311658059e-11 luc = 7.77352616871645e-18 wuc = 4.19664632264076e-17 puc = -1.01139651864783e-23
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0112296164664487 lu0 = -1.78583458343032e-09 wu0 = -6.52179043090389e-09 pu0 = 1.90552626059971e-15
+ a0 = 1.2288826280951 la0 = -1.47750595864118e-07 wa0 = -5.01094225701041e-07 pa0 = 1.79768718405565e-13
+ keta = 0.0314663465664558 lketa = -1.58650158704661e-08 wketa = 1.98582715547467e-07 pketa = -1.3103166624714e-13
+ a1 = 0.0
+ a2 = 0.787386106746973 la2 = 3.06943955640516e-09 wa2 = 8.89246955721644e-08 pa2 = -2.16387575711393e-14
+ ags = -0.0476830074917975 lags = 3.78246594706559e-07 wags = -2.04938984343482e-06 pags = 1.42804688530844e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.291202147720405+0*(0.0/sqrt(l*w*mult))} lvoff = 9.5721254686757e-09 wvoff = 4.99480350440181e-07 pvoff = -3.05202758095579e-13
+ nfactor = {0.610241922543693+0*(0.1/sqrt(l*w*mult))} lnfactor = 2.460197786771e-07 wnfactor = 3.48076392060329e-06 pnfactor = 1.85243067824195e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 1.99636279357148 leta0 = -7.43146007854966e-07 weta0 = -7.26866095849569e-06 peta0 = 3.58590665994235e-12
+ etab = 0.0135140434666189 letab = -6.7367502650702e-09 wetab = -6.16006018278115e-08 petab = 3.06643321931085e-14
+ dsub = 0.233059130242816 ldsub = 4.1879369638293e-08 wdsub = -3.37321844178465e-07 pdsub = 1.01720007264324e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.275271878875414 lpclm = 1.70660113063432e-07 wpclm = 1.42623942752934e-06 ppclm = -6.96997385168564e-13
+ pdiblc1 = -0.371270110801464 lpdiblc1 = 2.26435329200651e-07 wpdiblc1 = 2.60034727413468e-07 ppdiblc1 = -2.98226937062971e-13
+ pdiblc2 = -0.0175397966267037 lpdiblc2 = 8.86518352822473e-09 wpdiblc2 = 6.03900240334085e-08 ppdiblc2 = -2.97926936765937e-14
+ pdiblcb = -0.24812338325364 lpdiblcb = 1.14076436475842e-08 wpdiblcb = -8.66268209748202e-07 ppdiblcb = 4.27363026060758e-13
+ drout = 2.20347302615153 ldrout = -5.93718975775542e-07 wdrout = -4.83921417594755e-06 pdrout = 2.38736824313361e-12
+ pscbe1 = 800012145.528787 lpscbe1 = -0.00599185088026388 wpscbe1 = -0.0613317892493797 ppscbe1 = 3.0257302245304e-8
+ pscbe2 = 6.18965708313068e-08 lpscbe2 = -1.58769788319556e-14 wpscbe2 = -3.70062040175393e-13 ppscbe2 = 1.11032969845702e-19
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -6.80796803745295e-09 lalpha0 = 3.40796313566097e-15 walpha0 = -6.45731223359516e-15 palpha0 = 3.18563750269736e-21
+ alpha1 = 1.973352e-10 lalpha1 = -4.80191528976e-17
+ beta0 = 3.38890209240018 lbeta0 = 2.95565646187871e-06 wbeta0 = -5.3792309108046e-08 pbeta0 = 1.1069215210608e-13
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = -29739831.0699415 lbgidl = 262.976420462822 wbgidl = 3626.32854912971 pbgidl = -5.11040706563382e-6
+ cgidl = 461.556270432166 lcgidl = -7.97018473424639e-05 wcgidl = 0.000466845001557909 pcgidl = -2.30312379378575e-10
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.481728178967838 lkt1 = -1.3187823124365e-08 wkt1 = 1.57660814174172e-07 pkt1 = -7.77800707430581e-14
+ kt2 = 0.0187994330498334 lkt2 = -3.65008122459388e-08 wkt2 = -6.34108329535685e-08 pkt2 = 3.12829735076476e-14
+ at = 17492.6238288657 lat = 0.0335025071634901 wat = 0.323069608566668 pat = -1.95561320725403e-7
+ ute = -0.484655752365456 lute = -9.10354880599812e-09 wute = 7.5678242551706e-07 pute = 8.87205642102133e-14
+ ua1 = 8.99330330902921e-10 lua1 = -2.06763688339668e-16 wua1 = -9.34422304184432e-16 pua1 = 3.73173394356254e-22
+ ub1 = 3.00978003221546e-19 lub1 = 1.26672690666489e-26 wub1 = 9.28744143157988e-25 pub1 = -1.57953374432056e-31
+ uc1 = -4.52399672431535e-11 luc1 = 3.43165751198029e-17 wuc1 = 3.96612237151117e-16 puc1 = -1.95663887851658e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.24e-6
+ sbref = 1.24e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.16 pmos
* DC IV MOS Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.006443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.71750521473078+0*(0.007356/sqrt(l*w*mult))} lvth0 = -6.96923080167183e-08 wvth0 = -5.17398519924263e-07 pvth0 = 1.11877838725504e-13
+ k1 = 0.42695925292975 lk1 = 9.75479320609852e-08 wk1 = -6.46549873209486e-07 pk1 = 1.51752511924942e-13
+ k2 = 0.0286002974671029 lk2 = -3.30092478589708e-08 wk2 = 2.26240876049351e-07 pk2 = -4.60777099897629e-14
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 310339.438323621 lvsat = -0.0419676276536423 wvsat = -1.07114846853863 pvsat = 1.90530179530974e-7
+ ua = -1.72255887449559e-09 lua = -9.0430029489466e-17 wua = 1.14071420215235e-15 pua = -2.1627677639231e-22
+ ub = 1.40227758887013e-18 lub = 8.63723833621064e-26 wub = -5.62303154072208e-26 pub = 1.11777018891929e-31
+ uc = 1.54233088824656e-13 luc = -2.80030820768359e-20 wuc = -1.43398978647041e-18 puc = 4.47014248769406e-25
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0046405726924412 lu0 = -1.82469849550892e-10 wu0 = 7.55490937453325e-09 pu0 = -1.51986971665575e-15
+ a0 = 0.768832093875613 la0 = -3.58028189682179e-08 wa0 = 1.36304528141361e-06 pa0 = -2.73847260976699e-13
+ keta = -0.220551369452623 lketa = 4.54604711101845e-08 wketa = -4.52696345184815e-08 pketa = -7.16931230867929e-14
+ a1 = 0.0
+ a2 = 0.804864934722957 la2 = -1.18382348561454e-09 wa2 = 4.59669680178922e-07 pa2 = -1.11855100635378e-13
+ ags = 2.14244295756457 lags = -1.54694277378326e-07 wags = 1.32764637083813e-05 pags = -2.30131566628341e-12
+ b0 = 0.0
+ b1 = 1.31755895762121e-23 lb1 = -3.2061216162963e-30 wb1 = -9.28845098453027e-29 pb1 = 2.26023308567363e-35
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0965116424245087+0*(0.0/sqrt(l*w*mult))} lvoff = -3.78034727090172e-08 wvoff = -3.71184297167839e-07 pvoff = -9.33369640759381e-14
+ nfactor = {2.1045437171627+0*(0.1/sqrt(l*w*mult))} lnfactor = -1.17600631421899e-07 wnfactor = -1.05752118997927e-05 pnfactor = 3.60559611200772e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = -3.93148819350829 leta0 = 6.99325395639051e-07 weta0 = 2.47750551522521e-05 peta0 = -4.21154713101481e-12
+ etab = 0.101521044353953 letab = -2.81521978469925e-08 wetab = 1.59902358048617e-07 petab = -2.32357550573018e-14
+ dsub = 0.833221164896261 ldsub = -1.04162859550207e-07 wdsub = -6.04947606141277e-07 pdsub = 1.66843524928832e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.82744607231801 lpclm = -2.07042850820502e-07 wpclm = -5.05802082336134e-06 ppclm = 8.80869535762673e-13
+ pdiblc1 = 1.50803741944381 lpdiblc1 = -2.30871606594175e-07 wpdiblc1 = -3.5394486120025e-06 ppdiblc1 = 6.26331739783834e-13
+ pdiblc2 = 0.0556183270986758 lpdiblc2 = -8.93696798286167e-09 wpdiblc2 = -2.17658331770215e-07 ppdiblc2 = 3.78670371279485e-14
+ pdiblcb = -0.513855059808429 lpdiblcb = 7.60702583570734e-08 wpdiblcb = 3.093815034815e-06 ppdiblcb = -5.36275710504763e-13
+ drout = -3.41358717287403 ldrout = 7.7312521893494e-07 wdrout = 1.89744583258323e-05 pdrout = -3.40740319610449e-12
+ pscbe1 = 799956623.111479 lpscbe1 = 0.00751886310240479 wpscbe1 = 0.219042104465188 ppscbe1 = -3.79683203037551e-8
+ pscbe2 = -3.34073801295645e-08 lpscbe2 = 7.31409398696089e-15 wpscbe2 = 2.92552359326006e-13 ppscbe2 = -5.02062929001691e-20
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.47713144194748e-08 lalpha0 = -4.27647629884293e-15 walpha0 = 2.3061829405697e-14 palpha0 = -3.9974913855247e-21
+ alpha1 = -2.47625714285714e-10 lalpha1 = 6.02567460628571e-17
+ beta0 = 32.5574984252139 lbeta0 = -4.1421714325555e-06 wbeta0 = 2.36719272658651e-06 pbeta0 = -4.78425504509757e-13
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -1.35193009207452e-11 lagidl = 2.76235596474523e-17 wagidl = 5.73243204373986e-16 pagidl = -1.39491854865957e-22
+ bgidl = 1759526409.76291 lbgidl = -172.420048048964 wbgidl = 8427.5508730041 pbgidl = -0.00117343024491258
+ cgidl = -276.986680114878 lcgidl = 0.000100013717157753 wcgidl = -0.00166730357699253 pcgidl = 2.89007067428731e-10
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.53592367299 wkt1 = -1.619771821234e-7
+ kt2 = -0.131201028226 wkt2 = 6.51468666562244e-8
+ at = 540602.318962161 lat = -0.0937899598308556 wat = -2.34238766058088 pat = 4.53045720234424e-7
+ ute = -1.07196157535862 lute = 1.33810275549513e-07 wute = 3.8982069438669e-06 pute = -6.75707395236002e-13
+ ua1 = -1.60817226263034e-10 lua1 = 5.12104979259819e-17 wua1 = 2.08275628143746e-15 pua1 = -3.61020808311807e-22
+ ub1 = 2.54811740208192e-19 lub1 = 2.39012751757924e-26 wub1 = 9.72076683938877e-25 pub1 = -1.68497828240597e-31
+ uc1 = 9.57843492212001e-11 wuc1 = -4.07470511337231e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.17 pmos
* DC IV MOS Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.006443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.0161315323171252+0*(0.007356/sqrt(l*w*mult))} lvth0 = -1.91267019378936e-07 wvth0 = -4.89944538177174e-06 pvth0 = 8.71453077664422e-13
+ k1 = -0.392657687757268 lk1 = 2.39618693325791e-07 wk1 = 1.00916539780682e-06 pk1 = -1.35245861722483e-13
+ k2 = 0.803054948003311 lk2 = -1.67251668073616e-07 wk2 = -3.23722795959463e-06 pk2 = 5.54273051043092e-13
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 205485.824211048 lvsat = -0.0237925118905972 wvsat = -0.058712136199623 pvsat = 1.50364905559961e-8
+ ua = -6.21833455280008e-09 lua = 6.88858735036479e-16 wua = 3.7069846718057e-14 pua = -6.44416074843419e-21
+ ub = 4.43901906161463e-18 lub = -4.40010310040481e-25 wub = -2.68906774041579e-23 pub = 4.76320640836179e-30
+ uc = -5.68689044216977e-13 luc = 9.73067946203345e-20 wuc = 5.91137890799853e-18 puc = -8.2621726999245e-25
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = -0.0102124660880833 lu0 = 2.39212618658767e-09 wu0 = 1.14522258763292e-07 pu0 = -2.00613761250045e-14
+ a0 = 1.17101362378597 la0 = -1.05516160999819e-07 wa0 = -1.38328229199229e-05 pa0 = 2.36017414130656e-12
+ keta = 0.275607229049946 lketa = -4.05426680370539e-08 wketa = -2.58846860070149e-06 pketa = 3.69139899313439e-13
+ a1 = 0.0
+ a2 = -2.19600370085958 la2 = 5.18980744068992e-07 wa2 = 1.32486678338167e-05 pa2 = -2.32867446259064e-12
+ ags = 1.25
+ b0 = 0.0
+ b1 = -3.07430423444949e-23 lb1 = 4.40664620357521e-30 wb1 = 2.16730522972373e-28 pb1 = -3.1065719701814e-35
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {0.574511853609982+0*(0.0/sqrt(l*w*mult))} lvoff = -1.54117343464644e-07 wvoff = -6.80142001570368e-06 pvoff = 1.02126723490363e-12
+ nfactor = {-13.723479233335+0*(0.1/sqrt(l*w*mult))} lnfactor = 2.62599721077148e-06 wnfactor = 9.20303850035655e-05 pnfactor = -1.41798528440266e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = -1.51940007829828 leta0 = 2.81218865924778e-07 weta0 = 6.35996843866777e-06 peta0 = -1.01951283025552e-12
+ etab = -0.231132122977319 letab = 2.95092368718757e-08 wetab = -1.11565828990309e-07 petab = 2.38199975476516e-14
+ dsub = 0.0999383576860371 ldsub = 2.29429156859987e-08 wdsub = 2.06610389251714e-06 pdsub = -2.96151199745622e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 3.71862137087371 lpclm = -5.3485539472155e-07 wpclm = -1.12835390361757e-05 ppclm = 1.95998841173549e-12
+ pdiblc1 = 0.924450429477843 lpdiblc1 = -1.29713804927454e-07 wpdiblc1 = 4.27021779990339e-07 ppdiblc1 = -6.12083050234236e-14
+ pdiblc2 = 0.0339848896858175 lpdiblc2 = -5.18707120859164e-09 wpdiblc2 = -8.40619177647916e-08 ppdiblc2 = 1.47097019170764e-14
+ pdiblcb = -1.28618179332612 lpdiblcb = 2.09943829691563e-07 wpdiblcb = 6.11615581363059e-06 ppdiblcb = -1.0601622164231e-12
+ drout = 1.26942818544336 ldrout = -3.861929724508e-08 wdrout = -3.94695129404574e-06 pdrout = 5.65748104585929e-13
+ pscbe1 = 1037237333.48986 lpscbe1 = -41.1222449124662 wpscbe1 = -1197.98737433922 ppscbe1 = 0.000207656735493214
+ pscbe2 = 1.14644682539838e-08 lpscbe2 = -4.63902468146611e-16 wpscbe2 = -9.38564160314656e-15 ppscbe2 = 2.13103630488838e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 18.6713885325858 lbeta0 = -1.73518091598713e-06 wbeta0 = -2.95954589535218e-05 pbeta0 = 5.06191661241687e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 8.37890482199508e-10 lagidl = -1.19958109339046e-16 wagidl = -4.67218093371007e-15 pagidl = 7.69739474381258e-22
+ bgidl = -1130940033.82741 lbgidl = 328.607624350096 wbgidl = 13478.3817633864 pbgidl = -0.00204893116978967
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = 0.164051748335465 lkt1 = -1.21332339581714e-07 wkt1 = -6.8075615838838e-07 pkt1 = 8.9924110187821e-14
+ kt2 = -0.175354045021279 lkt2 = 7.65339562526016e-09 wkt2 = 3.76414252415214e-07 pkt2 = -5.39544661126921e-14
+ at = -184329.302219754 lat = 0.0318682375215751 wat = 1.56736426415516 pat = -2.24662858895472e-7
+ ute = -0.3
+ ua1 = 1.3462e-10
+ ub1 = 3.927e-19
+ uc1 = 3.71945786510145e-10 luc1 = -4.78692712167912e-17 wuc1 = -2.35433744980576e-15 puc1 = 3.37466021380258e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.18 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.004443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.0537489431687+0*(0.005856/sqrt(l*w*mult))} wvth0 = 5.86524686695862e-8
+ k1 = 0.44205207135451 wk1 = -5.80141215968923e-8
+ k2 = 0.0248237253676165 wk2 = -5.31710770688974e-9
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 323282.33637695 wvsat = -0.822955660079779
+ ua = -1.10744223691828e-09 wua = 2.78940299102583e-15
+ ub = 1.2393304653032e-18 wub = -8.11355992844838e-25
+ uc = -9.27767945288183e-12 wuc = -2.72434533704855e-16
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.00853738103508001 wu0 = 1.26067771702569e-8
+ a0 = 1.3101985775754 wa0 = -5.83783413380071e-7
+ keta = -0.012282397655245 wketa = 3.7473305957607e-8
+ a1 = 0.0
+ a2 = 1.07716489714687 wa2 = -8.45281483187463e-7
+ ags = 0.309122196092176 wags = -4.08481756909438e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.278390185468769+0*(0.0/sqrt(l*w*mult))} wvoff = -5.73912519381443e-8
+ nfactor = {1.41438576175584+0*(0.1/sqrt(l*w*mult))} wnfactor = 1.51744570432627e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.347005573953947 wpclm = -6.04564498173483e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 0.000133338415931977 wpdiblc2 = 1.78567236809097e-10
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 865373846.835292 wpscbe1 = -330.121073140511
+ pscbe2 = 7.8629967022153e-09 wpscbe2 = 6.13072686726336e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.25320264185616e-10 walpha0 = -6.32835026573253e-16
+ alpha1 = 2.5248701384693e-10 walpha1 = -7.70020108774829e-16
+ beta0 = 1.27556883885757 wbeta0 = 2.56304465703625e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 1831914799.42999 wbgidl = -1461.96803056708
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.423448049072474 wkt1 = -6.36549844626647e-8
+ kt2 = -0.0472892886219128 wkt2 = -1.63933688432524e-8
+ at = 90000.0
+ ute = -0.154755494649972 wute = -5.0278340702204e-8
+ ua1 = 1.72985419276207e-09 wua1 = 1.15892950575362e-15
+ ub1 = -7.7370399143252e-19 wub1 = 1.07442513567083e-25
+ uc1 = 1.1396316068919e-10 wuc1 = -1.02636045017316e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.19 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.004443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.0537489431687+0*(0.005856/sqrt(l*w*mult))} wvth0 = 5.86524686695879e-8
+ k1 = 0.44205207135451 wk1 = -5.80141215968931e-8
+ k2 = 0.0248237253676165 wk2 = -5.3171077068898e-9
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 323282.33637695 wvsat = -0.822955660079779
+ ua = -1.10744223691828e-09 wua = 2.78940299102583e-15
+ ub = 1.2393304653032e-18 wub = -8.11355992844838e-25
+ uc = -9.2776794528818e-12 wuc = -2.72434533704855e-16
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.00853738103508001 wu0 = 1.26067771702568e-8
+ a0 = 1.3101985775754 wa0 = -5.83783413380071e-7
+ keta = -0.012282397655245 wketa = 3.7473305957607e-8
+ a1 = 0.0
+ a2 = 1.07716489714687 wa2 = -8.45281483187465e-7
+ ags = 0.309122196092176 wags = -4.08481756909438e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.278390185468769+0*(0.0/sqrt(l*w*mult))} wvoff = -5.73912519381438e-8
+ nfactor = {1.41438576175584+0*(0.1/sqrt(l*w*mult))} wnfactor = 1.51744570432627e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.347005573953947 wpclm = -6.04564498173483e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 0.000133338415931977 wpdiblc2 = 1.78567236809097e-10
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 865373846.835292 wpscbe1 = -330.12107314051
+ pscbe2 = 7.8629967022153e-09 wpscbe2 = 6.13072686726336e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.25320264185616e-10 walpha0 = -6.32835026573253e-16
+ alpha1 = 2.5248701384693e-10 walpha1 = -7.70020108774829e-16
+ beta0 = 1.27556883885757 wbeta0 = 2.56304465703625e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 1831914799.42999 wbgidl = -1461.96803056707
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.423448049072474 wkt1 = -6.36549844626656e-8
+ kt2 = -0.0472892886219128 wkt2 = -1.63933688432524e-8
+ at = 90000.0
+ ute = -0.154755494649972 wute = -5.02783407022042e-8
+ ua1 = 1.72985419276207e-09 wua1 = 1.15892950575362e-15
+ ub1 = -7.7370399143252e-19 wub1 = 1.07442513567083e-25
+ uc1 = 1.1396316068919e-10 wuc1 = -1.02636045017318e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.20 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.004443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.06262269978816+0*(0.005856/sqrt(l*w*mult))} lvth0 = 7.09309359890674e-08 wvth0 = 6.99529191074277e-08 pvth0 = -9.03283199018835e-14
+ k1 = 0.530793050435021 lk1 = -7.09336640241456e-07 wk1 = -4.27339440244663e-07 pk1 = 2.95214210390933e-12
+ k2 = -0.00610486988431966 lk2 = 2.47222715713921e-07 wk2 = 1.25899871399314e-07 pk2 = -1.04886166533482e-12
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 548343.001603383 lvsat = -1.79898596765972 wvsat = -1.43743032144168 pvsat = 4.91170366070124e-6
+ ua = -1.64119992627694e-09 lua = 4.26650562114275e-15 wua = 4.70334052511315e-15 pua = -1.52987496208464e-20
+ ub = 1.44675049405168e-18 lub = -1.65797839775631e-24 wub = -1.40676265850699e-24 pub = 4.75928672609059e-30
+ uc = 5.95594457962296e-12 luc = -1.21767505856734e-16 wuc = -3.59605785576392e-16 puc = 6.96789280092326e-22
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.00587205428747613 lu0 = 2.13048575740384e-08 wu0 = 2.25511735555569e-08 pu0 = -7.94889215136818e-14
+ a0 = 1.32862577376842 la0 = -1.47294807563097e-07 wa0 = -6.15368556722904e-07 pa0 = 2.52470726517685e-13
+ keta = -0.0129741666777652 lketa = 5.52954361493362e-09 wketa = 6.91001360601783e-08 pketa = -2.52803942878427e-13
+ a1 = 0.0
+ a2 = 1.35386817615754 la2 = -2.21178283484059e-06 wa2 = -1.68915515006468e-06 pa2 = 6.74536744864898e-12
+ ags = 0.348472695282173 lags = -3.14541840494371e-07 wags = -1.0100218765759e-06 pags = 4.8083134970545e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.277638024913813+0*(0.0/sqrt(l*w*mult))} lvoff = -6.01227354603256e-09 wvoff = -6.61957634316593e-08 pvoff = 7.03774362925567e-14
+ nfactor = {1.4504189948289+0*(0.1/sqrt(l*w*mult))} lnfactor = -2.8802581118571e-07 wnfactor = 1.67945572669866e-06 pnfactor = -1.29500086821006e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.212075360148291 lpclm = 1.07854280536088e-06 wpclm = -9.96685515937816e-07 ppclm = 3.13435583189431e-12
+ pdiblc1 = 0.39
+ pdiblc2 = 0.000322784426404387 lpdiblc2 = -1.51430599445751e-09 wpdiblc2 = -4.69556414514648e-10 ppdiblc2 = 5.18067141082484e-15
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 930638813.52868 lpscbe1 = -521.684938338991 wpscbe1 = -659.692329633705 ppscbe1 = 0.00263437444823481
+ pscbe2 = 6.3331713917849e-09 lpscbe2 = 1.22284107872252e-14 wpscbe2 = 1.18984913767618e-14 ppscbe2 = -4.61036912288251e-20
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.20364460368239e-10 lalpha0 = 3.96134149739854e-17 walpha0 = -6.07809494901723e-16 palpha0 = -2.00037533280245e-22
+ alpha1 = 2.53834796508647e-10 lalpha1 = -1.0773282365639e-17 walpha1 = -7.76826063758127e-16 palpha1 = 5.44022985942843e-23
+ beta0 = -9.69692649132035 lbeta0 = 8.77068638775337e-05 wbeta0 = 7.94311761784672e-05 pbeta0 = -4.30047416404189e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.54406130953349e-10 lagidl = -4.34886593982381e-16 wagidl = -2.74736935413853e-16 pagidl = 2.1960651858471e-21
+ bgidl = 1435802806.08597 lbgidl = 3166.25704865253 wbgidl = 819.438396469894 pbgidl = -0.0182360526866788
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.368870747285083 lkt1 = -4.36254820314618e-07 wkt1 = -2.04077764051027e-07 pkt1 = 1.12244674014928e-12
+ kt2 = -0.0431578686030913 lkt2 = -3.30238366304066e-08 wkt2 = -3.27594345306962e-08 pkt2 = 1.30819494769942e-13
+ at = 12613.5593365334 lat = 0.618575976840033 wat = 0.368994300011135 pat = -2.9494961600624e-6
+ ute = -0.027887934724782 lute = -1.0140952877173e-06 wute = -4.84842005339567e-07 pute = 3.47361425396509e-12
+ ua1 = 1.27911773946639e-09 lua1 = 3.60288882011355e-15 wua1 = 2.31592881441541e-15 pua1 = -9.24828653990001e-21
+ ub1 = -6.24466392744989e-19 lub1 = -1.19290656861779e-24 wub1 = 2.14706081627819e-25 pub1 = -8.57393954595471e-31
+ uc1 = 3.57861121649557e-10 luc1 = -1.94955883946702e-15 wuc1 = -2.05101149701663e-17 puc1 = 8.19038214947304e-23
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.21 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.004443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.05461346271302+0*(0.005856/sqrt(l*w*mult))} lvth0 = 3.89473452259103e-08 wvth0 = 5.27721241651509e-08 pvth0 = -2.17195985887146e-14
+ k1 = 0.373015378371156 lk1 = -7.92770668372826e-08 wk1 = 7.58194485716647e-08 pk1 = 9.42858593161316e-13
+ k2 = 0.0458286860643386 lk2 = 3.98344732690177e-08 wk2 = -4.14704549886032e-08 pk2 = -3.8049538089755e-13
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 98301.1165003386 lvsat = -0.00181660628610292 wvsat = -0.193012368399835 pvsat = -5.76778390629876e-8
+ ua = 1.15223286153522e-10 lua = -2.74748593713789e-15 wua = 3.35712147503249e-16 pua = 2.14266674934153e-21
+ ub = 6.77593851070971e-19 lub = 1.41352405261099e-24 wub = 1.60576913336901e-25 pub = -1.49962994505735e-30
+ uc = -6.04314185481519e-11 luc = 1.43339674041208e-16 wuc = -1.38651508798689e-16 puc = -1.85555829626594e-22
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0143527239856468 lu0 = -1.25613229971153e-08 wu0 = 5.68288302050885e-10 pu0 = 8.29616951878358e-15
+ a0 = 1.03422763702158 la0 = 1.02833645903724e-06 wa0 = 7.48612711297419e-07 pa0 = -5.19436750235606e-12
+ keta = -0.0141123846217396 lketa = 1.00748325828883e-08 wketa = 5.02574710229668e-08 pketa = -1.77558812564059e-13
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.332223406673803 lags = -2.496529388216e-07 wags = -7.72526473189937e-07 pags = 3.85991407788799e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.275784622900298+0*(0.0/sqrt(l*w*mult))} lvoff = -1.34135342358804e-08 wvoff = -5.92838911275679e-08 pvoff = 4.27759939694741e-14
+ nfactor = {1.63005129719678+0*(0.1/sqrt(l*w*mult))} lnfactor = -1.00535831025887e-06 wnfactor = 7.94968055319523e-07 pnfactor = 2.23705736043976e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.280058625165649 leta0 = -7.98901710101742e-07 weta0 = -6.1012723164166e-07 peta0 = 2.43644425894945e-12
+ etab = -0.244894021371516 letab = 6.98410941515688e-07 wetab = 5.33381677504415e-07 petab = -2.12997332128213e-12
+ dsub = 1.31493822630977 ldsub = -3.0147235067754e-06 wdsub = -2.30236696717005e-06 pdsub = 9.19412949994492e-12
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.0135958562374929 lpclm = 1.97972424926045e-06 wpclm = 1.29082362683677e-06 ppclm = -6.00044135329489e-12
+ pdiblc1 = 0.39
+ pdiblc2 = -0.000867982236533001 lpdiblc2 = 3.24082776978356e-09 wpdiblc2 = 3.30281662860508e-09 ppdiblc2 = -9.88368921244079e-15
+ pdiblcb = 0.0109618223819394 lpdiblcb = -1.43607711867049e-07 wpdiblcb = -1.81597932070984e-07 ppdiblcb = 7.2518192286048e-13
+ drout = 0.56
+ pscbe1 = 829062731.07521 lpscbe1 = -116.057308386416 wpscbe1 = -88.6338374073166 ppscbe1 = 0.000353944871004461
+ pscbe2 = 8.69514328830249e-09 lpscbe2 = 2.79625865792938e-15 wpscbe2 = 3.94168111007434e-15 ppscbe2 = -1.4329458432072e-20
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.84803028897529e-10 lalpha0 = -2.17711569399633e-16 walpha0 = -9.33207653711671e-16 palpha0 = 1.09938729942555e-21
+ alpha1 = 4.01770528127303e-10 lalpha1 = -6.01530660996222e-16 walpha1 = -1.52386337060073e-15 palpha1 = 3.03757476342652e-21
+ beta0 = 13.6788228296188 lbeta0 = -5.64040416424703e-06 wbeta0 = -4.32571733337314e-05 pbeta0 = 5.9888631860156e-11
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 8.07229865515796e-11 lagidl = -1.40644893483307e-16 wagidl = 9.73439483004568e-17 pagidl = 7.10220453837163e-22
+ bgidl = 2584536810.133 lbgidl = -1421.02610160067 wbgidl = -4832.42877731601 pbgidl = 0.00433376326935304
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.505091761503496 lkt1 = 1.07721732162309e-07 wkt1 = 2.25418313307938e-07 pkt1 = -5.92676266419217e-13
+ kt2 = -0.0753600598698912 lkt2 = 9.55703974385738e-08 wkt2 = 8.74969746462684e-08 pkt2 = -3.4940499373998e-13
+ at = 175682.251731657 lat = -0.0326124291117261 wat = -0.336473176143857 pat = -1.32326079768581e-7
+ ute = -1.41237058533168 lute = 4.51461189129194e-06 wute = 6.54266887837163e-06 pute = -2.45896120033724e-11
+ ua1 = 3.14777222840417e-10 lua1 = 7.4538264500957e-15 wua1 = 1.28574877453173e-14 pua1 = -5.13442943979099e-20
+ ub1 = 4.71851051745124e-19 lub1 = -5.57087267976306e-24 wub1 = -8.92903366267034e-24 pub1 = 3.56566494284207e-29
+ uc1 = -5.31956518410092e-10 luc1 = 1.6037837556535e-15 wuc1 = 7.97928326735067e-16 puc1 = -3.18639750842756e-21
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.22 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.004443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.02932531166733+0*(0.005856/sqrt(l*w*mult))} lvth0 = -1.14604872032017e-08 wvth0 = -5.11874586806516e-08 pvth0 = 1.85506988361975e-13
+ k1 = 0.10039887683441 lk1 = 4.6413976510297e-07 wk1 = 1.35716335838934e-06 pk1 = -1.61129291334682e-12
+ k2 = 0.162272482600208 lk2 = -1.92277371230199e-07 wk2 = -5.64890412770687e-07 pk2 = 6.62857510907873e-13
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 244068.671580339 lvsat = -0.292380612994161 wvsat = -0.834859689580168 pvsat = 1.22174081644397e-6
+ ua = -1.73563971923514e-09 lua = 9.41909624297528e-16 wua = 4.54063758214276e-15 pua = -6.2391709066919e-21
+ ub = 1.62637248106967e-18 lub = -4.77712444153367e-25 wub = -2.23604560110502e-24 pub = 3.27764878463528e-30
+ uc = 5.31004707896902e-11 luc = -8.2967755187707e-17 wuc = -4.62924689993097e-16 puc = 4.60830224829106e-22
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.00595722128274793 lu0 = 4.17375156967585e-09 wu0 = 1.87828087659224e-08 pu0 = -2.80115262736291e-14
+ a0 = 3.05232777324131 la0 = -2.99441923029471e-06 wa0 = -6.79709899743419e-06 pa0 = 9.84678638370358e-12
+ keta = 0.10088003799562 lketa = -2.19143933132354e-07 wketa = -4.16135307794606e-07 pketa = 7.52119636378603e-13
+ a1 = 0.0
+ a2 = 0.8
+ ags = -1.64763899562792 lags = 3.69688202245772e-06 wags = 6.67208527632395e-06 pags = -1.09797134176645e-11
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.313009896080735+0*(0.0/sqrt(l*w*mult))} lvoff = 6.07890173550665e-08 wvoff = 8.76984374480882e-08 pvoff = -2.50209466908865e-13
+ nfactor = {0.214745534570712+0*(0.1/sqrt(l*w*mult))} lnfactor = 1.81582444800265e-06 wnfactor = 5.22948181832324e-06 pnfactor = -6.60242743487854e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = -0.727385830331298 leta0 = 1.20927560592963e-06 weta0 = 1.22025446328332e-06 peta0 = -1.21212512804893e-12
+ etab = -34.2820315755331 letab = 6.8545930639453e-05 wetab = 0.000173116659082056 petab = -3.46146778336317e-10
+ dsub = -0.65187505261954 ldsub = 9.0580014101899e-07 wdsub = 4.60473393434011e-06 pdsub = -4.57405719686954e-12
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.8471449765229 lpclm = -1.72936116083248e-06 wpclm = -5.0051780124959e-06 ppclm = 6.54961796244923e-12
+ pdiblc1 = 0.390866386212638 lpdiblc1 = -1.72700056032672e-09 wpdiblc1 = 3.94632362357761e-08 ppdiblc1 = -7.86635683917507e-14
+ pdiblc2 = 0.00108351045437734 lpdiblc2 = -6.49156767730276e-10 wpdiblc2 = -3.30005931961042e-09 ppdiblc2 = 3.27807432442317e-15
+ pdiblcb = -0.121021474460452 lpdiblcb = 1.19479609094169e-07 wpdiblcb = 3.6330656746386e-07 ppdiblcb = -3.60996922433307e-13
+ drout = 0.230293343769541 ldrout = 6.57216806717111e-07 wdrout = 4.01420155559661e-07 pdrout = -8.00166050042983e-13
+ pscbe1 = 741874537.849581 lpscbe1 = 57.7382303215727 wpscbe1 = 177.267674814635 ppscbe1 = -0.00017608671756502
+ pscbe2 = 1.32054628524648e-08 lpscbe2 = -6.19433272145884e-15 wpscbe2 = -7.67765136125417e-15 ppscbe2 = 8.83179851766105e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.5066333061691e-10 lalpha0 = -1.4965961150834e-16 walpha0 = -7.6081097860876e-16 palpha0 = 7.55742455869269e-22
+ alpha1 = 1.0e-10
+ beta0 = 12.673999595604 lbeta0 = -3.63745182860242e-06 wbeta0 = -2.59283534049786e-05 pbeta0 = 2.53464366010158e-11
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -7.90704969165552e-11 lagidl = 1.77877529266097e-16 wagidl = 9.04259845054499e-16 pagidl = -8.98235665966746e-22
+ bgidl = 2578052665.42636 lbgidl = -1408.10100955941 wbgidl = -5413.76045930138 pbgidl = 0.00549255380165839
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.391249452887838 lkt1 = -1.19204467609008e-07 wkt1 = -3.30145970616336e-07 pkt1 = 5.14751132169828e-13
+ kt2 = -0.0110141705813727 lkt2 = -3.26927088240231e-08 wkt2 = -1.56002906015875e-07 pkt2 = 1.35972571379336e-13
+ at = 351979.590328345 lat = -0.384032613435371 wat = -1.10422113114352 pat = 1.39805509335454e-6
+ ute = 1.6847753734155 lute = -1.65904683982524e-06 wute = -1.02711048508271e-05 pute = 8.92592209444106e-12
+ ua1 = 3.686021553228e-09 lua1 = 7.33797019049587e-16 wua1 = -1.30744886405701e-14 pua1 = 3.46899547182051e-22
+ ub1 = -7.5076055188382e-19 lub1 = -3.13379451100854e-24 wub1 = 4.47378850369363e-24 pub1 = 8.94029469696506e-30
+ uc1 = 7.14555127546979e-10 luc1 = -8.80935275675275e-16 wuc1 = -2.40395057058658e-15 puc1 = 3.19602936900178e-21
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.23 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.004443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.08326102983466+0*(0.005856/sqrt(l*w*mult))} lvth0 = 4.21159112097006e-08 wvth0 = 1.95472327421469e-07 pvth0 = -5.9509550245132e-14
+ k1 = 0.606367207056303 lk1 = -3.84578041029854e-08 wk1 = -2.92454366424754e-07 pk1 = 2.73350581845565e-14
+ k2 = -0.0564653548022676 lk2 = 2.50032346995016e-08 wk2 = 1.26709642120851e-07 pk2 = -2.41351044179779e-14
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -131455.051406357 lvsat = 0.080641370949998 wvsat = 0.613173136561131 pvsat = -2.16645215009572e-7
+ ua = -1.85246834309527e-11 lua = -7.63765991138129e-16 wua = -4.56847092988074e-15 pua = 2.80925272442449e-21
+ ub = 8.33963468675203e-19 lub = 3.0941753940053e-25 wub = 2.26089752279267e-24 pub = -1.189335704171e-30
+ uc = -4.1567900070096e-11 luc = 1.10699349854114e-17 wuc = -3.40471374250269e-17 puc = 3.48098545162443e-23
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0138438141188205 lu0 = -3.66030078492281e-09 wu0 = -2.19898639878834e-08 pu0 = 1.24895189342909e-14
+ a0 = -0.66051158659657 la0 = 6.93685193727924e-07 wa0 = 5.40905712830643e-06 pa0 = -2.27805232992735e-12
+ keta = -0.221735743270409 lketa = 1.01322581798881e-07 wketa = 6.65604950141895e-07 pketa = -3.22414067959525e-13
+ a1 = 0.0
+ a2 = 0.855668795604156 la2 = -5.52979300878407e-08 wa2 = -2.93726959638508e-07 pa2 = 2.91770150633396e-13
+ ags = 3.4206042760025 lags = -1.33759661249711e-06 wags = -9.58669614967402e-06 pags = 5.17075200647346e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.27415565940833+0*(0.0/sqrt(l*w*mult))} lvoff = 2.21936276073727e-08 wvoff = 3.79378951534595e-09 pvoff = -1.66863791740651e-13
+ nfactor = {2.2574641838547+0*(0.1/sqrt(l*w*mult))} lnfactor = -2.13285609639805e-07 wnfactor = -3.0519707134829e-06 pnfactor = 1.62385406016071e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.49
+ etab = 68.9839487907733 letab = -3.40320917656531e-05 wetab = -0.000348363542547731 petab = 1.71859322190214e-10
+ dsub = 0.224453312887367 ldsub = 3.53098750830884e-08 wdsub = 2.01607097438947e-08 pdsub = -2.00263990955808e-14
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.406119044464942 lpclm = 5.08891615247537e-07 wpclm = 3.16328859371136e-06 ppclm = -1.56443031922749e-12
+ pdiblc1 = 1.00904408541858 lpdiblc1 = -6.15786399934154e-07 wpdiblc1 = -1.36768834766852e-06 ppdiblc1 = 1.31911357166057e-12
+ pdiblc2 = 0.000666837698516518 lpdiblc2 = -2.35259885769001e-10 wpdiblc2 = -1.19596932074974e-09 ppdiblc2 = 1.1880017731349e-15
+ pdiblcb = 0.220530859393146 lpdiblcb = -2.19797303111296e-07 wpdiblcb = -2.21406643782003e-10 ppdiblcb = 1.09228310830117e-16
+ drout = 0.785275872460918 ldrout = 1.05931571631876e-07 wdrout = -8.02840311119321e-07 pdrout = 3.96071633406984e-13
+ pscbe1 = 800000000.0
+ pscbe2 = 2.53824092974694e-08 lpscbe2 = -1.82901563492468e-14 wpscbe2 = -6.0826192132795e-14 ppscbe2 = 6.16262637105818e-20
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.57425481733679 lbeta0 = 4.3498044995201e-07 wbeta0 = -6.08391403110394e-07 pbeta0 = 1.95156186004012e-13
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 2.6182827825113e-10 lagidl = -1.60750178261421e-16 wagidl = -8.17191085838074e-16 pagidl = 8.11746958824222e-22
+ bgidl = 772337411.716175 lbgidl = 385.584569130557 wbgidl = 1896.52550630667 pbgidl = -0.00176903103884678
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.514009554323414 lkt1 = 2.73780603080502e-09 wkt1 = 3.73609188019475e-07 pkt1 = -1.84315609599152e-13
+ kt2 = -0.0328143309139654 lkt2 = -1.10377811595661e-08 wkt2 = -3.79820865533236e-08 pkt2 = 1.87380066160436e-14
+ at = -134217.756003195 lat = 0.0989256861749088 wat = 0.579587741575663 pat = -2.7453624465459e-7
+ ute = 0.342407017985139 lute = -3.25621342378752e-07 wute = -2.55351331173964e-06 pute = 1.25974515018701e-12
+ ua1 = 8.51884992919061e-09 lua1 = -4.06683505427237e-15 wua1 = -2.61261316584609e-14 pua1 = 1.33115925192877e-20
+ ub1 = -8.24516964542902e-18 lub1 = 4.31068682915546e-24 wub1 = 2.69950423496756e-23 pub1 = -1.3430922555895e-29
+ uc1 = -3.66276989096027e-10 luc1 = 1.92696337406656e-16 wuc1 = 1.61618783423289e-15 puc1 = -7.97326873764784e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.24 pmos
* DC IV MOS Parameters
+ lmin = 2.5e-07 lmax = 5e-07 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.006443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.951832437393914+0*(0.007356/sqrt(l*w*mult))} lvth0 = -2.27228077278341e-08 wvth0 = 7.7280948571156e-10 pvth0 = 3.65431205342582e-14
+ k1 = 0.163421034192796 lk1 = 1.80064374925152e-07 wk1 = -7.40544611169513e-08 pk1 = -8.04099143001847e-14
+ k2 = 0.113533628240646 lk2 = -5.88637235969233e-08 wk2 = 1.28297159411033e-08 pk2 = 3.20461906036865e-14
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 25456.3242167981 lvsat = 0.00323102672282168 wvsat = 0.136624734824863 pvsat = 1.84542204061952e-8
+ ua = -9.29658715624296e-10 lua = -3.1426894996393e-16 wua = 1.3525292982704e-15 pua = -1.11801686131143e-22
+ ub = 1.02857980744732e-18 lub = 2.13405904063373e-25 wub = 4.09831504818267e-26 pub = -9.41675875639128e-32
+ uc = -4.75896127117167e-11 luc = 1.40406746566033e-17 wuc = 1.21163496857495e-16 puc = -4.17614493794266e-23
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.00899873800679532 lu0 = -1.27004062596853e-09 wu0 = 4.74357066987863e-09 pu0 = -6.99100252900136e-16
+ a0 = 0.571238059801894 la0 = 8.60162866729989e-08 wa0 = 2.81984130340993e-06 pa0 = -1.00069377330456e-12
+ keta = 0.101631076408027 lketa = -5.8206558287639e-08 wketa = -1.55731081685113e-07 pketa = 8.27822073099479e-14
+ a1 = 0.0
+ a2 = 0.688662408791688 la2 = 2.70926667694481e-08 wa2 = 5.87453919277015e-07 pa2 = -1.4294986180903e-13
+ ags = -2.81930579041722 lags = 1.74078813985027e-06 wags = 1.19465906859851e-05 pags = -5.45243665445695e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0860307542340639+0*(0.0/sqrt(l*w*mult))} lvoff = -7.06155368614891e-08 wvoff = -5.36582293480602e-07 pvoff = 9.97242642924044e-14
+ nfactor = {1.58868573574939+0*(0.1/sqrt(l*w*mult))} lnfactor = 1.16648212391568e-07 wnfactor = -1.46012509327047e-06 pnfactor = 8.38536125576345e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.366482927314561 leta0 = 6.09356656044893e-08 weta0 = 9.61812183072228e-07 peta0 = -4.74498498772486e-13
+ etab = 0.00464865828736444 letab = -1.98179689275993e-09 wetab = -1.68326921688757e-08 petab = 6.65304348992104e-15
+ dsub = 0.294072112845111 ldsub = 9.6427554953515e-10 wdsub = -6.45421677173141e-07 pdsub = 3.08330684501296e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.794166853835649 lpclm = -8.32550292482797e-08 wpclm = -1.19404642489531e-06 ppclm = 5.85208624181893e-13
+ pdiblc1 = -0.801818314507566 lpdiblc1 = 2.77580834720609e-07 wpdiblc1 = 2.43419216080237e-06 ppdiblc1 = -5.56498554627437e-13
+ pdiblc2 = -0.0043274684194413 lpdiblc2 = 2.22862110585207e-09 wpdiblc2 = -6.32882727505457e-09 ppdiblc2 = 3.72023565059574e-15
+ pdiblcb = -0.567731063497013 lpdiblcb = 1.6908225740349e-07 wpdiblcb = 7.47668180620868e-07 ppdiblcb = -3.68853124891138e-13
+ drout = 1.00440263087424 ldrout = -2.17198511023697e-09 wdrout = 1.21578219985483e-06 pdrout = -5.99791558911982e-13
+ pscbe1 = 800000000.0
+ pscbe2 = -4.3110488492554e-08 lpscbe2 = 1.54999928606878e-14 wpscbe2 = 1.60196538590211e-13 ppscbe2 = -4.74126482188446e-20
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -2.05703849742862e-08 lalpha0 = 1.01974863824444e-14 walpha0 = 6.30393453463266e-14 palpha0 = -3.10997045544661e-20
+ alpha1 = 3.4575883349272e-10 lalpha1 = -1.21242171397631e-16 walpha1 = -7.49501085525521e-16 palpha1 = 3.6975736653099e-22
+ beta0 = -6.47112278601071 lbeta0 = 7.85743694603227e-06 wbeta0 = 4.97367914124534e-05 pbeta0 = -2.46420356138606e-11
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 3.43185516096839e-09 lagidl = -1.72464490052739e-15 wagidl = -1.68250096106299e-14 pagidl = 8.70901213420795e-21
+ bgidl = 213203934.577475 lbgidl = 661.42636047521 wbgidl = 2399.52516351304 pbgidl = -0.00201717988373366
+ cgidl = 586.270015136891 lcgidl = -0.000141227876727604 wcgidl = -0.000162927257997569 pcgidl = 8.03782076060047e-11
+ egidl = 1.97886865382484 legidl = -9.26917303940642e-07 wegidl = -9.48780232947651e-06 pegidl = 4.68069342561929e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.400324591436112 lkt1 = -5.33473061900915e-08 wkt1 = -2.53406317016177e-07 pkt1 = 1.25014965624127e-13
+ kt2 = 0.0915056319202278 lkt2 = -7.23695429842614e-08 wkt2 = -4.30558393590991e-07 pkt2 = 2.12410816777392e-13
+ at = 66816.0075095094 lat = -0.000251908648921745 wat = 0.0739992365477296 pat = -2.51102227611195e-8
+ ute = -0.33479019576 lute = 8.46577665584692e-9
+ ua1 = 4.29498206488999e-10 lua1 = -7.60504540981951e-17 wua1 = 1.4381088013842e-15 pua1 = -2.86894740691394e-22
+ ub1 = 5.51281263333473e-19 lub1 = -2.89366692716141e-26 wub1 = -3.35222792226797e-25 pub1 = 5.21357886808695e-32
+ uc1 = 1.17907496082509e-11 luc1 = 6.18115532976476e-18 wuc1 = 1.08621819570329e-16 puc1 = -5.35872712231869e-23
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.24e-6
+ sbref = 1.24e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.25 pmos
* DC IV MOS Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.006443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.872075470773442+0*(0.007356/sqrt(l*w*mult))} lvth0 = -4.21307084713266e-08 wvth0 = 2.63141424879187e-07 pvth0 = -2.73011335983598e-14
+ k1 = 0.5872654990847 lk1 = 7.69269105272855e-08 wk1 = -1.45605508934173e-06 pk1 = 2.55883354570775e-13
+ k2 = -0.0286485264068586 lk2 = -2.42654024493088e-08 wk2 = 5.15332677866063e-07 pk2 = -9.02318751452093e-14
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -56002.2210168059 lvsat = 0.0230529862028764 wvsat = 0.778782468250751 pvsat = -1.37807158130194e-7
+ ua = -1.94484830035453e-09 lua = -6.72347467948452e-17 wua = 2.26321849652601e-15 pua = -3.3340697425626e-22
+ ub = 1.74686672431862e-18 lub = 3.8619402285744e-26 wub = -1.79631661434303e-24 pub = 3.52917262609037e-31
+ uc = 3.47284410300679e-11 luc = -5.99043590481514e-18 wuc = -1.76024826658942e-16 puc = 3.05557628884162e-23
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.00513970925320032 lu0 = -3.30992287126226e-10 wu0 = 5.034398420105e-09 pu0 = -7.69869695984721e-16
+ a0 = 3.33141756518768 la0 = -5.85640273808568e-07 wa0 = -1.15773507141778e-05 pa0 = 2.50269013787121e-12
+ keta = -0.0806582499923219 lketa = -1.3848638180031e-08 wketa = -7.51693823346802e-07 pketa = 2.2780258894042e-13
+ a1 = 0.0
+ a2 = 0.558328548562314 la2 = 5.88078476499434e-08 wa2 = 1.7046148732098e-06 pa2 = -4.14797574017127e-13
+ ags = 11.9724486774532 lags = -1.85860780885238e-06 wags = -3.63625310015815e-05 pags = 6.30300839875213e-12
+ b0 = 0.0
+ b1 = -1.31755895762121e-23 lb1 = 3.2061216162963e-30 wb1 = 4.01821515404542e-29 pb1 = -9.77784439155104e-36
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0961063178566346+0*(0.0/sqrt(l*w*mult))} lvoff = -6.81637693607001e-08 wvoff = -3.73231081742935e-07 pvoff = 5.99747071305837e-14
+ nfactor = {-2.06280383418596+0*(0.1/sqrt(l*w*mult))} lnfactor = 1.0051943813605e-06 wnfactor = 1.04688188923193e-05 pnfactor = -2.06422924598909e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 1.59573856023088 leta0 = -2.38188941598102e-07 weta0 = -3.13601503507358e-06 peta0 = 5.22658580836678e-13
+ etab = 0.0406813692995357 letab = -1.07499247250397e-08 wetab = 4.67127032605198e-07 petab = -1.11112748017153e-13
+ dsub = 0.166883633834733 ldsub = 3.19140656549622e-08 wdsub = 2.75988514390392e-06 pdsub = -5.20309866725955e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.0335155624375654 lpclm = 1.18151554562812e-07 wpclm = 4.33935567624487e-06 ppclm = -7.61278376305355e-13
+ pdiblc1 = 0.66815501043113 lpdiblc1 = -8.01195342233238e-08 wpdiblc1 = 7.01741031826505e-07 ppdiblc1 = -1.34927361804708e-13
+ pdiblc2 = 0.00562324910435547 lpdiblc2 = -1.92766594953582e-10 wpdiblc2 = 3.48039233699959e-08 ppdiblc2 = -6.28892562586955e-15
+ pdiblcb = 0.910068479288695 lpdiblcb = -1.90522527738899e-07 wpdiblcb = -4.0966317501371e-06 ppdiblcb = 8.09949131659644e-13
+ drout = 1.53850669319406 ldrout = -1.32139799427018e-07 wdrout = -6.03233904801292e-06 pdrout = 1.16395176930166e-12
+ pscbe1 = 800000000.0
+ pscbe2 = 4.8803272583498e-08 lpscbe2 = -6.86611793203657e-15 wpscbe2 = -1.2259024296869e-13 ppscbe2 = 2.14001216321354e-20
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 7.39228034795937e-08 lalpha0 = -1.27962971095458e-14 walpha0 = -2.25140519094024e-13 palpha0 = 3.90254072987199e-20
+ alpha1 = -7.77710119616857e-10 lalpha1 = 1.52140516714147e-16 walpha1 = 2.67678959116258e-15 palpha1 = -4.63989354152939e-22
+ beta0 = 68.4900003161139 lbeta0 = -1.03834528273925e-05 wbeta0 = -0.000179082678423471 pbeta0 = 3.10384365370736e-11
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -1.21942749144563e-08 lagidl = 2.0777863397663e-15 wagidl = 6.20829188539313e-14 pagidl = -1.04922853625014e-20
+ bgidl = 7131481718.19918 lbgidl = -1022.05351883573 wbgidl = -18699.4385445206 pbgidl = 0.00311699974705182
+ cgidl = -722.392911203183 lcgidl = 0.000177219542442137 wcgidl = 0.000581883064277032 pcgidl = -1.00862446595652e-10
+ egidl = -6.61024519223159 legidl = 1.16314048113104e-06 wegidl = 3.3885008319559e-05 pegidl = -5.87355957209572e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.860500726041802 lkt1 = 5.86310340525878e-08 wkt1 = 1.47705325982393e-06 pkt1 = -2.96071606884989e-13
+ kt2 = -0.436632348495648 lkt2 = 5.6146496894177e-08 wkt2 = 1.60749629382358e-06 pkt2 = -2.83525334748695e-13
+ at = 153765.342308894 lat = -0.0214099858803345 wat = -0.38896065505447 pat = 8.75455113415765e-8
+ ute = -0.3
+ ua1 = 7.32574130346422e-11 lua1 = 1.06364680994012e-17 wua1 = 9.00739697426206e-16 pua1 = -1.56132417672464e-22
+ ub1 = 5.30588259791808e-19 lub1 = -2.39012751757925e-26 wub1 = -4.20523644771641e-25 pub1 = 7.28927275374267e-32
+ uc1 = 3.7192270660305e-11 wuc1 = -1.11595619642564e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.26 pmos
* DC IV MOS Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.006443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.58932328220464+0*(0.007356/sqrt(l*w*mult))} lvth0 = 8.21955926665348e-08 wvth0 = 3.04476738632712e-06 pvth0 = -5.09462614503821e-13
+ k1 = -0.0350215001207808 lk1 = 1.84792894395565e-07 wk1 = -7.96805151148258e-07 pk1 = 1.41610288784197e-13
+ k2 = -0.159538280445407 lk2 = -1.57723426377513e-09 wk2 = 1.62361968753711e-06 pk2 = -2.82340128827568e-13
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 169619.735154785 lvsat = -0.0160558724359948 wvsat = 0.122402367256745 pvsat = -2.40315441840944e-8
+ ua = 6.45831239663715e-09 lua = -1.52382181568999e-15 wua = -2.69439523370175e-14 pua = 4.7293056036885e-21
+ ub = -5.18513091974681e-18 lub = 1.24019800991276e-24 wub = 2.17087988958522e-23 pub = -3.72141244969719e-30
+ uc = 7.31852179223179e-13 luc = -9.7535186587409e-20 wuc = -6.56018990846856e-19 puc = 1.576845048439e-25
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0285603820110996 lu0 = -4.39068486163497e-09 wu0 = -8.12706284973415e-08 pu0 = 1.41900710598316e-14
+ a0 = -5.61744441828076 la0 = 9.65537564681884e-07 wa0 = 2.04471401280309e-05 pa0 = -3.04837105573556e-12
+ keta = -0.705107081218503 lketa = 9.43920733270528e-08 wketa = 2.36388583800499e-06 pketa = -3.12245758398976e-13
+ a1 = 0.0
+ a2 = 2.44215683986062 la2 = -2.67731180707122e-07 wa2 = -1.01728471790329e-05 pa2 = 1.64401794319453e-12
+ ags = 1.25
+ b0 = 0.0
+ b1 = 3.07430423444949e-23 lb1 = -4.40664620357521e-30 wb1 = -9.3758353594393e-29 pb1 = 1.34391348875131e-35
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.980044083558183+0*(0.0/sqrt(l*w*mult))} lvoff = 8.50562350704748e-08 wvoff = 1.04868670247494e-06 pvoff = -1.86497677750175e-13
+ nfactor = {15.3361089942057+0*(0.1/sqrt(l*w*mult))} lnfactor = -2.01069837048726e-06 wnfactor = -5.47130439836701e-05 pnfactor = 9.23426450120916e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.149907636831496 leta0 = 1.24284990021005e-08 weta0 = -2.06960517520864e-06 peta0 = 3.37809228547409e-13
+ etab = -0.0502303205623976 letab = 5.00852577224816e-09 wetab = -1.025073294701e-06 petab = 1.47542272317449e-13
+ dsub = 0.785782032553578 ldsub = -7.53645449821647e-08 wdsub = -1.39722985506456e-06 pdsub = 2.00276132965244e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.41917561129315 lpclm = -1.33655028109323e-07 wpclm = 3.28069252589311e-07 ppclm = -6.59700102017489e-14
+ pdiblc1 = 1.09673359026096 lpdiblc1 = -1.54408488093867e-07 wpdiblc1 = -4.42963767365563e-07 ppdiblc1 = 6.34934786776462e-14
+ pdiblc2 = 0.0114313462497088 lpdiblc2 = -1.19953053793484e-09 wpdiblc2 = 2.98276622840598e-08 ppdiblc2 = -5.42635048175556e-15
+ pdiblcb = -0.188015344889178 lpdiblcb = -1.82873823554952e-10 wpdiblcb = 5.70698356334438e-07 ppdiblcb = 9.23465664080792e-16
+ drout = -0.293204208071499 ldrout = 1.85365304776552e-07 wdrout = 3.94393944657323e-06 pdrout = -5.65316392392914e-13
+ pscbe1 = 800000000.0
+ pscbe2 = 1.03975245252142e-08 lpscbe2 = -2.08942375109786e-16 wpscbe2 = -3.99785083095377e-15 ppscbe2 = 8.43553563764412e-22
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 10.5299447529672 lbeta0 = -3.36772716187804e-07 wbeta0 = 1.15167332693456e-05 pbeta0 = -1.99968428693587e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -8.98817400935598e-10 lagidl = 1.19854325287652e-16 wagidl = 4.09774615282994e-15 pagidl = -4.41251496837919e-22
+ bgidl = 2358841974.44934 lbgidl = -194.773690933619 wbgidl = -4144.11771260946 pbgidl = 0.000594009544690016
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = 0.278988308483013 lkt1 = -1.38885716213875e-07 wkt1 = -1.26115615648829e-06 pkt1 = 1.78564136919738e-13
+ kt2 = -0.0685659549787205 lkt2 = -7.65339562526016e-09 wkt2 = -1.62838072330096e-07 pkt2 = 2.33408836116513e-14
+ at = -6781.76583984483 lat = 0.00641892875195169 wat = 0.670794977191492 pat = -9.61504104406741e-8
+ ute = -0.3
+ ua1 = 1.3462e-10
+ ub1 = 3.927e-19
+ uc1 = 3.34046627238648e-11 luc1 = 6.56536384486661e-19 wuc1 = -6.44792050586758e-16 puc1 = 9.24232029470047e-23
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.27 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 2e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.004443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.034517+0*(0.005856/sqrt(l*w*mult))}
+ k1 = 0.42302944
+ k2 = 0.023080264
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 53438.0
+ ua = -1.9280657e-10
+ ub = 9.7328962e-19
+ uc = -9.8608028e-11
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0126711
+ a0 = 1.118778
+ keta = 4.9707517e-6
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.17518243
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.29720858+0*(0.0/sqrt(l*w*mult))}
+ nfactor = {1.911951+0*(0.1/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.14877095
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00019189
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 757128280.0
+ pscbe2 = 9.873241e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.7815831e-11
+ alpha1 = 6.3056523e-17
+ beta0 = 9.6797043
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 1352540500.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.4443203
+ kt2 = -0.052664618
+ at = 90000.0
+ ute = -0.17124159
+ ua1 = 2.1098632e-9
+ ub1 = -7.3847396e-19
+ uc1 = 1.1059776e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.28 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 2e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.004443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.034517+0*(0.005856/sqrt(l*w*mult))}
+ k1 = 0.42302944
+ k2 = 0.023080264
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 53438.0
+ ua = -1.9280657e-10
+ ub = 9.7328962e-19
+ uc = -9.8608028e-11
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0126711
+ a0 = 1.118778
+ keta = 4.9707517e-6
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.17518243
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.29720858+0*(0.0/sqrt(l*w*mult))}
+ nfactor = {1.911951+0*(0.1/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.14877095
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00019189
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 757128280.0
+ pscbe2 = 9.873241e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.7815831e-11
+ alpha1 = 6.3056523e-17
+ beta0 = 9.6797043
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 1352540500.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.4443203
+ kt2 = -0.052664618
+ at = 90000.0
+ ute = -0.17124159
+ ua1 = 2.1098632e-9
+ ub1 = -7.3847396e-19
+ uc1 = 1.1059776e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.29 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 2e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.004443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.0396853777065+0*(0.005856/sqrt(l*w*mult))} lvth0 = 4.13125899197166e-8
+ k1 = 0.390669914700905 lk1 = 2.58660623235218e-7
+ k2 = 0.0351772658317135 lk2 = -9.66954244275052e-8
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 77014.5327768425 lvsat = -0.188455195353381
+ ua = -9.89907109822351e-11 lua = -7.49901870889343e-16
+ ub = 9.85477846643321e-19 lub = -9.74246151806612e-26
+ uc = -1.11957558265434e-10 luc = 1.06707307552848e-16
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0132665066958 lu0 = -4.75928696699256e-9
+ a0 = 1.126848536098 la0 = -6.45105228725166e-8
+ keta = 0.00968353076963815 lketa = -7.73640015766657e-08 wketa = -2.99852972050473e-24 pketa = 4.18096279767136e-29
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.017289988568175 lags = 1.26208765200978e-6
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.299343388544765+0*(0.0/sqrt(l*w*mult))} lvoff = 1.70642462635953e-8
+ nfactor = {2.00110676335525+0*(0.1/sqrt(l*w*mult))} lnfactor = -7.12652151146524e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.114734399685775 lpclm = 2.10628732484659e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 0.000168818489705 lpdiblc2 = 1.84418379958414e-10
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 714327962.84966 lpscbe1 = 342.117401489868
+ pscbe2 = 1.02346458760091e-08 lpscbe2 = -2.88883132878883e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.1065813124638e-11 lalpha0 = -2.59782056161896e-17
+ alpha1 = -8.83803561262884e-13 lalpha1 = 7.06504462287938e-18 walpha1 = 2.34440593327997e-34 palpha1 = -2.72457263015603e-39
+ beta0 = 16.3482835524884 lbeta0 = -5.33042079449267e-05 wbeta0 = 1.35525271560688e-20
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 6.43208327881951e-11 lagidl = 2.85195643082475e-16
+ bgidl = 1704493843.79725 lbgidl = -2813.28203720162
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.435787145678045 lkt1 = -6.82083867015476e-8
+ kt2 = -0.0538995747481865 lkt2 = 9.87142670363557e-9
+ at = 133605.523841315 lat = -0.348553690730689
+ ute = -0.18686596419218 lute = 1.24890903956571e-7
+ ua1 = 2.0385028489407e-09 lua1 = 5.70407405815647e-16
+ ub1 = -5.54065005497301e-19 lub1 = -1.47404310356671e-24
+ uc1 = 3.51135925346025e-10 luc1 = -1.92270285751067e-15 puc1 = -7.52316384526264e-37
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.30 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 2e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.004443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.0373096643247+0*(0.005856/sqrt(l*w*mult))} lvth0 = 3.1825563395068e-8
+ k1 = 0.39787631532893 lk1 = 2.29883029764101e-7
+ k2 = 0.0322306662092167 lk2 = -8.4928656184203e-08 pk2 = 5.04870979341448e-29
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 35013.023362553 lvsat = -0.0207289717519407
+ ua = 2.2530214708257e-10 lua = -2.04491286412814e-15
+ ub = 7.3024646981917e-19 lub = 9.21800540683538e-25
+ uc = -1.05894772401041e-10 luc = 8.24965543747024e-17
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0145390637694 lu0 = -9.84103748616824e-9
+ a0 = 1.279695175654 la0 = -6.74878816783792e-7
+ keta = 0.00236686763209579 lketa = -4.81460926363186e-8
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.0789146275940702 lags = 1.01599963925139e-6
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.29522360732579+0*(0.0/sqrt(l*w*mult))} lvoff = 6.12567370175419e-10
+ nfactor = {1.8907185940324+0*(0.1/sqrt(l*w*mult))} lnfactor = -2.71834879839156e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.40966078061423 lpclm = 1.22001243377312e-8
+ pdiblc1 = 0.39
+ pdiblc2 = 0.000215
+ pdiblcb = -0.0485835162604495 lpdiblcb = 9.41769516564709e-8
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 9.9876069955871e-09 lpscbe2 = -1.90232158012222e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -2.1192557782444e-11 lalpha0 = 1.42773752745155e-16
+ alpha1 = -9.78990408614235e-11 lalpha1 = 3.94479678312628e-16 walpha1 = -2.00296714216273e-32 palpha1 = 5.87747175411144e-38
+ beta0 = -0.5050558384638 lbeta0 = 1.39968726718593e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.1264173309365e-10 lagidl = 9.223395569849e-17
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.43117787025461 lkt1 = -8.66147814024163e-8
+ kt2 = -0.046670102192069 lkt2 = -1.89983007746655e-8
+ at = 65353.85212337 lat = -0.0760016964958941
+ ute = 0.73294808402065 lute = -3.54823748770556e-06 pute = 8.07793566946316e-28
+ ua1 = 4.5307033248294e-09 lua1 = -9.38179145816879e-15
+ ub1 = -2.45594843985464e-18 lub1 = 6.12082028642297e-24
+ uc1 = -2.7031855873761e-10 luc1 = 5.5897494905091e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.31 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 2e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.004443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.0461095036822+0*(0.005856/sqrt(l*w*mult))} lvth0 = 4.93666175802695e-8
+ k1 = 0.5454080839698 lk1 = -6.41976508749532e-8
+ k2 = -0.0229531449202714 lk2 = 2.50713315250285e-08 wk2 = -2.64697796016969e-23
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -29678.9552125639 lvsat = 0.108224007437026
+ ua = -2.46780240508461e-10 lua = -1.10389310181221e-15
+ ub = 8.93180803063241e-19 lub = 5.97017342723469e-25
+ uc = -9.86909462006041e-11 luc = 6.81368938639756e-17 wuc = 9.86076131526265e-32
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0121160398104 lu0 = -5.01113175378311e-9
+ a0 = 0.823582341108001 la0 = 2.34308228604462e-7
+ keta = -0.0355693011631478 lketa = 2.74735141976547e-8
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.540114866427681 lags = 9.6671677575281e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.28425387944166+0*(0.0/sqrt(l*w*mult))} lvoff = -2.12538080709204e-8
+ nfactor = {1.9294746740774+0*(0.1/sqrt(l*w*mult))} lnfactor = -3.49088846923895e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = -0.32726858 leta0 = 8.1182393672004e-07 peta0 = -2.01948391736579e-28
+ etab = 22.482326763364 letab = -4.49544099258305e-05 wetab = 6.67038445962762e-21 petab = 1.81753552562921e-26
+ dsub = 0.858001400000001 ldsub = -5.940175146732e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.20596428508744 lpclm = 4.18236089338113e-7
+ pdiblc1 = 0.40380624592792 lpdiblc1 = -2.75205146454682e-8
+ pdiblc2 = 1.43233000000041e-06 lpdiblc2 = 4.2571255218246e-10
+ pdiblcb = -0.00189449793638372 lpdiblcb = 1.10995724841425e-9
+ drout = 0.361917635016081 ldrout = 3.94845105252317e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 1.06879873224826e-08 lpscbe2 = -3.29841630017542e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.19602200021408e-12 lalpha0 = 9.81457458983515e-17
+ alpha1 = 1.0e-10
+ beta0 = 4.17218150587221 lbeta0 = 4.67355773837533e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 2.1743320265992e-10 lagidl = -1.166508626638e-16
+ bgidl = 802899192.027401 lbgidl = 392.888530362486
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.499503183520001 lkt1 = 4.95806618913891e-8
+ kt2 = -0.0621669880280001 lkt2 = 1.18922306437575e-8
+ at = -10090.7286459999 lat = 0.0743848532457603
+ ute = -1.6830846545 lute = 1.26773237923172e-06 pute = 1.61558713389263e-27
+ ua1 = -6.0105839752e-10 lua1 = 8.47544189935722e-16 wua1 = 3.94430452610506e-31
+ ub1 = 7.16179343460001e-19 lub1 = -2.02302564913869e-25
+ uc1 = -7.3692013666e-11 luc1 = 1.67031784950957e-16 wuc1 = 2.46519032881566e-32 puc1 = -4.70197740328915e-38
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.32 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 2e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.004443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.0191663245768+0*(0.005856/sqrt(l*w*mult))} lvth0 = 2.26029339340693e-8
+ k1 = 0.510472424072761 lk1 = -2.94947323441472e-8
+ k2 = -0.014917698045952 lk2 = 1.70894167977859e-08 wk2 = 6.61744490042422e-24
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 69602.315528176 lvsat = 0.0096041485219607
+ ua = -1.5165106213508e-09 lua = 1.57378335232961e-16
+ ub = 1.5753040065058e-18 lub = -8.05615559377584e-26
+ uc = -5.27318395745652e-11 luc = 2.24839668062795e-17 puc = 2.35098870164458e-38
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0066334131912 lu0 = 4.34969606879774e-10
+ a0 = 1.113099680712 la0 = -5.32803464830964e-8
+ keta = -0.00348616462015639 lketa = -4.39588448968728e-9
+ a1 = 0.0
+ a2 = 0.75935673367364 la2 = 4.03725008860937e-8
+ ags = 0.27715951215524 lags = 3.57875223277559e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.27291168884736+0*(0.0/sqrt(l*w*mult))} lvoff = -3.25204369914811e-8
+ nfactor = {1.2567334619324+0*(0.1/sqrt(l*w*mult))} lnfactor = 3.19170563265793e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.49
+ etab = -45.243261151015 letab = 2.2319990121863e-5
+ dsub = 0.23106394041644 ldsub = 2.87432875546143e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.63111242831704 lpclm = -4.07971696129197e-9
+ pdiblc1 = 0.5605837704226 lpdiblc1 = -1.83253587271965e-7
+ pdiblc2 = 0.00027468346307008 lpdiblc2 = 1.54281818160893e-10
+ pdiblcb = 0.220458260914565 lpdiblcb = -2.1976148752307e-07 wpdiblcb = -1.65436122510606e-23 ppdiblcb = -2.60324098722934e-29
+ drout = 0.52202728996784 ldrout = 2.35802100821846e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 5.43770966587601e-09 lpscbe2 = 1.91688400668287e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.3747653643888 lbeta0 = 4.98971493524154e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -6.12587401724004e-12 lagidl = 1.05418863444537e-16
+ bgidl = 1394201615.9452 lbgidl = -194.474636807173
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.39150438388 lkt1 = -5.76986497454087e-8
+ kt2 = -0.045268526732 lkt2 = -4.89365310308857e-9
+ at = 55827.075188 lat = 0.00890619382090246
+ ute = -0.494881232720001 lute = 8.74447686476191e-8
+ ua1 = -4.78189710399998e-11 lua1 = 2.97990444514932e-16
+ ub1 = 6.0641208816e-19 lub1 = -9.32665790686782e-26
+ uc1 = 1.6366545464e-10 luc1 = -6.87444079011883e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.33 pmos
* DC IV MOS Parameters
+ lmin = 2.5e-07 lmax = 5e-07 wmin = 2e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.006443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.951579035816+0*(0.007356/sqrt(l*w*mult))} lvth0 = -1.07404439286061e-8
+ k1 = 0.1391388305636 lk1 = 1.53698240010475e-7
+ k2 = 0.117740448063352 lk2 = -4.8355887687486e-08 pk2 = 1.26217744835362e-29
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 70255.10584 lvsat = 0.00928210225510609
+ ua = -4.861690008968e-10 lua = -3.50928339118574e-16
+ ub = 1.0420180418272e-18 lub = 1.82528675304853e-25
+ uc = -7.860517951676e-12 luc = 3.47238739486535e-19
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.01055413854848 lu0 = -1.49927319943003e-9
+ a0 = 1.49585434488 la0 = -2.42107766994409e-7
+ keta = 0.050567389226496 lketa = -3.10625566372871e-08 pketa = 6.31088724176809e-30
+ a1 = 0.0
+ a2 = 0.88128653265272 la2 = -1.97801022826473e-8
+ ags = 1.097940292214 lags = -4.70471251950703e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.26197424659896+0*(0.0/sqrt(l*w*mult))} lvoff = -3.79162928754222e-8
+ nfactor = {1.1099157291336+0*(0.1/sqrt(l*w*mult))} lnfactor = 3.91601329929288e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.68185784099488 leta0 = -9.4650763560732e-8
+ etab = -0.000870723701341264 letab = 1.99713232889716e-10
+ dsub = 0.0824405601279197 ldsub = 1.02064848739392e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.402643129340079 lpclm = 1.08632870057404e-7
+ pdiblc1 = -0.00365505965856028 lpdiblc1 = 9.51068686826147e-8
+ pdiblc2 = -0.00640266916101696 lpdiblc2 = 3.44847360702274e-09 wpdiblc2 = -8.27180612553028e-25 ppdiblc2 = -1.18329135783152e-30
+ pdiblcb = -0.3225732332316 lpdiblcb = 4.8136583736011e-8
+ drout = 1.40305344137712 ldrout = -1.98841578662106e-07 wdrout = -1.6940658945086e-21
+ pscbe1 = 800000000.0
+ pscbe2 = 9.4174066817368e-09 lpscbe2 = -4.64517597278701e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 9.8374004106232 lbeta0 = -2.22601954915029e-07 wbeta0 = 1.35525271560688e-20
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -2.08500774325672e-09 lagidl = 1.1310102870514e-15 pagidl = 1.88079096131566e-37
+ bgidl = 1000000000.0
+ cgidl = 532.846726441352 lcgidl = -0.000114872138329124
+ egidl = -1.1321491658048 legidl = 6.07866005159808e-07 wegidl = 4.2351647362715e-22
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.48341565304 lkt1 = -1.23553280405526e-8
+ kt2 = -0.049672987568 lkt2 = -2.72076520317801e-9
+ at = 91080.103192 lat = -0.00848546450853489 wat = 1.11022302462516e-16
+ ute = -0.33479019576 lute = 8.46577665584692e-9
+ ua1 = 9.01049146559999e-10 lua1 = -1.70122254885617e-16 wua1 = -7.88860905221012e-31 pua1 = -1.88079096131566e-37
+ ub1 = 4.4136286032e-19 lub1 = -1.18415231045482e-26
+ uc1 = 4.74074714316e-11 luc1 = -1.13899269811227e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.24e-6
+ sbref = 1.24e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.34 pmos
* DC IV MOS Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 2e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.006443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.785792300714286+0*(0.007356/sqrt(l*w*mult))} lvth0 = -5.10826564747872e-8
+ k1 = 0.109830032788 lk1 = 1.60830184243594e-7
+ k2 = 0.140327289931343 lk2 = -5.38521246139591e-8
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 199357.877371429 lvsat = -0.0221335079638087
+ ua = -1.20274672320286e-09 lua = -1.76557749328064e-16
+ ub = 1.15786067182571e-18 lub = 1.54339761406275e-25
+ uc = -2.29894954758249e-11 luc = 4.02869387225787e-18
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.00679047121599999 lu0 = -5.83429918079006e-10
+ a0 = -0.464755998 la0 = 2.34983232621324e-7
+ keta = -0.327136074690686 lketa = 6.08470488653921e-8
+ a1 = 0.0
+ a2 = 1.117265914878 la2 = -7.72028531945827e-8
+ ags = 0.0492995661671429 lags = 2.0812701179972e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.218487508549715+0*(0.0/sqrt(l*w*mult))} lvoff = -4.84982687388495e-8
+ nfactor = {1.36988594933714+0*(0.1/sqrt(l*w*mult))} lnfactor = 3.28340696485398e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.567449993717428 leta0 = -6.68109868199316e-8
+ etab = 0.193850720008982 letab = -4.71834134366929e-08 wetab = 5.02512222125964e-23 petab = 7.34626717987067e-30
+ dsub = 1.07184049999343 ldsub = -1.38693753827601e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.38934427018857 lpclm = -1.31469012154387e-7
+ pdiblc1 = 0.898253486238858 lpdiblc1 = -1.24361753058971e-7
+ pdiblc2 = 0.0170353361227257 lpdiblc2 = -2.25488372271263e-9
+ pdiblcb = -0.433203011048126 lpdiblcb = 7.50570126103288e-8
+ drout = -0.439476576346856 ldrout = 2.49515990790811e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 8.60635267050002e-09 lpscbe2 = 1.50908501258472e-16
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 9.76940471184571 lbeta0 = -2.06056017565912e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 8.16250109563771e-09 lagidl = -1.36259801878749e-15
+ bgidl = 1000000000.0
+ cgidl = -531.595451576257 lcgidl = 0.000144147092385325 wcgidl = -2.16840434497101e-19 pcgidl = -2.58493941422821e-26
+ egidl = 4.50053273501714 legidl = -7.62779543222401e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.376180031714286 lkt1 = -3.84498296627092e-8
+ kt2 = 0.0904601689714285 lkt2 = -3.68204872491695e-8
+ at = 26226.4785142858 lat = 0.00729588681329076
+ ute = -0.3
+ ua1 = 3.68606868285714e-10 lua1 = -4.05588157749091e-17
+ ub1 = 3.927e-19
+ uc1 = 6.0045e-13
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.35 pmos
* DC IV MOS Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 2e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.006443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {0.563947705288165+0*(0.007356/sqrt(l*w*mult))} lvth0 = -2.85043889635241e-07 wvth0 = -3.52215401226537e-06 pvth0 = 6.10523132178055e-13
+ k1 = 1.1621400030665 lk1 = -2.15751213845409e-08 wk1 = -4.44783910763394e-06 pk1 = 7.70979535239053e-13
+ k2 = 0.196801235004252 lk2 = -6.3641205305007e-08 wk2 = 5.36876029742731e-07 pk2 = -9.30610172435454e-14
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 166575.3705211 lvsat = -0.0164510537913863 wvsat = 0.131686894552284 pvsat = -2.28263429279037e-8
+ ua = -9.19908293852142e-09 lua = 1.20951117756283e-15 wua = 2.08070669586988e-14 pua = -3.60665537248692e-21
+ ub = 6.49203981318285e-18 lub = -7.70276182598288e-25 wub = -1.39035614649683e-23 pub = 2.41001553721467e-30
+ uc = -3.94304914786051e-13 luc = 1.12088730788524e-19 wuc = 2.77846982258246e-18 puc = -4.81614402106797e-25
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = -0.0202401630908956 lu0 = 4.10200617140966e-09 wu0 = 6.75584532832165e-08 pu0 = -1.17104471752062e-14
+ a0 = -1.65176677274049 la0 = 4.40737306293291e-07 wa0 = 8.35284566083008e-06 pa0 = -1.44786556115696e-12
+ keta = -0.450576214903672 lketa = 8.22439158896306e-08 wketa = 1.58763231380209e-06 pketa = -2.75197010009826e-13
+ a1 = 0.0
+ a2 = -0.893484834715332 la2 = 2.71336660238426e-7
+ ags = -10.3645163606705 lags = 2.0132370369259e-06 wags = 3.54212806777271e-05 pags = -6.13985395011586e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {0.296966117646507+0*(0.0/sqrt(l*w*mult))} lvoff = -1.3784596939645e-07 wvoff = -2.84586519796949e-06 pvoff = 4.93296581685636e-13
+ nfactor = {-16.1671722290247+0*(0.1/sqrt(l*w*mult))} lnfactor = 3.36817928700628e-06 wnfactor = 4.13638422012832e-05 pnfactor = -7.16992567948602e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = -1.01574925099338 leta0 = 2.0761760385975e-07 weta0 = 1.48534782631153e-06 peta0 = -2.57467221517188e-13
+ etab = -0.250295517592581 letab = 2.98040070966869e-08 wetab = -4.14926020566733e-07 petab = 7.19224465529963e-14
+ dsub = 0.330562837006492 ldsub = -1.02021662807714e-08 wdsub = -8.92866415455878e-09 pdsub = 1.54767678722307e-15
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.43122109036495 lpclm = -3.12065856410121e-07 wpclm = -2.75840855325518e-06 ppclm = 4.78137021804147e-13
+ pdiblc1 = 0.95148729129 lpdiblc1 = -1.33589194358926e-7
+ pdiblc2 = 0.0212117343376133 lpdiblc2 = -2.97881223648482e-9
+ pdiblcb = -0.245247273470374 lpdiblcb = 4.24771409700764e-08 wpdiblcb = 7.45240984115895e-07 ppdiblcb = -1.29178581704681e-13
+ drout = 1.0
+ pscbe1 = 617872337.420839 lpscbe1 = 31.5696447761463 wpscbe1 = 555.442418355022 ppscbe1 = -9.62792779128233e-5
+ pscbe2 = 6.53942374298324e-09 lpscbe2 = 5.09185827696371e-16 wpscbe2 = 7.76836193646916e-15 ppscbe2 = -1.34655232134369e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 14.9251119737245 lbeta0 = -1.09973600292546e-06 wbeta0 = -1.88739367985472e-06 pbeta0 = 3.27157045678659e-13
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -7.68430126385546e-10 lagidl = 1.85471737375578e-16 wagidl = 3.70009857929166e-15 pagidl = -6.41367687537257e-22
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.279092992818759 lkt1 = -5.5278702810782e-08 wkt1 = 4.40847939122636e-07 pkt1 = -7.64157000716393e-14
+ kt2 = -0.102764678099045 lkt2 = -3.3272787076678e-09 wkt2 = -5.85407832439275e-08 pkt2 = 1.01473422859359e-14
+ at = 94560.1438756112 lat = -0.00454893407311069 wat = 0.361728278503676 pat = -6.27012563392702e-8
+ ute = 0.55761956064625 lute = -1.486580594033e-07 wute = -2.61551856564833e-06 pute = 4.5336875713235e-13
+ ua1 = 1.39125024527775e-10 lua1 = -7.80891941595511e-19 wua1 = -1.37391634143906e-17 pua1 = 2.38151910792368e-24
+ ub1 = 3.04264409813457e-19 lub1 = 1.53292483317552e-26 wub1 = 2.69705751373809e-25 pub1 = -4.67502555316328e-32
+ uc1 = -4.86875125689353e-10 luc1 = 8.4498041338841e-17 wuc1 = 9.41927175944102e-16 puc1 = -1.63271772823799e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.36 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.004443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.034517+0*(0.005856/sqrt(l*w*mult))}
+ k1 = 0.42302944
+ k2 = 0.023080264
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 53438.0
+ ua = -1.9280657e-10
+ ub = 9.7328962e-19
+ uc = -9.8608028e-11
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0126711
+ a0 = 1.118778
+ keta = 4.9707517e-6
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.17518243
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.29720858+0*(0.0/sqrt(l*w*mult))}
+ nfactor = {1.911951+0*(0.1/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.14877095
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00019189
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 757128280.0
+ pscbe2 = 9.873241e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.7815831e-11
+ alpha1 = 6.3056523e-17
+ beta0 = 9.6797043
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 1352540500.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.4443203
+ kt2 = -0.052664618
+ at = 90000.0
+ ute = -0.17124159
+ ua1 = 2.1098632e-9
+ ub1 = -7.3847396e-19
+ uc1 = 1.1059776e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.37 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.004443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.034517+0*(0.005856/sqrt(l*w*mult))}
+ k1 = 0.42302944
+ k2 = 0.023080264
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 53438.0
+ ua = -1.9280657e-10
+ ub = 9.7328962e-19
+ uc = -9.8608028e-11
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0126711
+ a0 = 1.118778
+ keta = 4.9707517e-6
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.17518243
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.29720858+0*(0.0/sqrt(l*w*mult))}
+ nfactor = {1.911951+0*(0.1/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.14877095
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00019189
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 757128280.0
+ pscbe2 = 9.873241e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.7815831e-11
+ alpha1 = 6.3056523e-17
+ beta0 = 9.6797043
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 1352540500.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.4443203
+ kt2 = -0.052664618
+ at = 90000.0
+ ute = -0.17124159
+ ua1 = 2.1098632e-9
+ ub1 = -7.3847396e-19
+ uc1 = 1.1059776e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.38 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.004443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.0396853777065+0*(0.005856/sqrt(l*w*mult))} lvth0 = 4.13125899197166e-8
+ k1 = 0.390669914700905 lk1 = 2.58660623235217e-7
+ k2 = 0.0351772658317135 lk2 = -9.66954244275053e-8
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 77014.5327768425 lvsat = -0.18845519535338
+ ua = -9.89907109822347e-11 lua = -7.49901870889345e-16
+ ub = 9.8547784664332e-19 lub = -9.74246151806642e-26
+ uc = -1.11957558265435e-10 luc = 1.06707307552848e-16
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0132665066958 lu0 = -4.75928696699256e-9
+ a0 = 1.126848536098 la0 = -6.45105228725098e-8
+ keta = 0.00968353076963815 lketa = -7.73640015766658e-08 wketa = -5.98413474393831e-24 pketa = 3.44140569902666e-29
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.0172899885681752 lags = 1.26208765200978e-6
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.299343388544765+0*(0.0/sqrt(l*w*mult))} lvoff = 1.70642462635944e-8
+ nfactor = {2.00110676335525+0*(0.1/sqrt(l*w*mult))} lnfactor = -7.12652151146537e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.114734399685775 lpclm = 2.1062873248466e-06 ppclm = 1.61558713389263e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 0.000168818489705 lpdiblc2 = 1.84418379958414e-10
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 714327962.849661 lpscbe1 = 342.117401489864
+ pscbe2 = 1.02346458760091e-08 lpscbe2 = -2.88883132878889e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.1065813124638e-11 lalpha0 = -2.59782056161897e-17 walpha0 = 4.93038065763132e-32
+ alpha1 = -8.83803561262885e-13 lalpha1 = 7.06504462287938e-18 walpha1 = -5.98843842082906e-34 palpha1 = -5.57183174346062e-39
+ beta0 = 16.3482835524884 lbeta0 = -5.33042079449269e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 6.43208327881949e-11 lagidl = 2.85195643082476e-16
+ bgidl = 1704493843.79725 lbgidl = -2813.28203720161
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.435787145678044 lkt1 = -6.82083867015476e-8
+ kt2 = -0.0538995747481865 lkt2 = 9.87142670363578e-9
+ at = 133605.523841315 lat = -0.348553690730689
+ ute = -0.18686596419218 lute = 1.2489090395657e-7
+ ua1 = 2.0385028489407e-09 lua1 = 5.70407405815647e-16
+ ub1 = -5.54065005497301e-19 lub1 = -1.4740431035667e-24
+ uc1 = 3.51135925346025e-10 luc1 = -1.92270285751067e-15 wuc1 = 3.94430452610506e-31
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.39 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.004443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.0373096643247+0*(0.005856/sqrt(l*w*mult))} lvth0 = 3.18255633950646e-8
+ k1 = 0.397876315328929 lk1 = 2.29883029764102e-7
+ k2 = 0.0322306662092167 lk2 = -8.49286561842029e-8
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 35013.0233625529 lvsat = -0.0207289717519407
+ ua = 2.25302147082569e-10 lua = -2.04491286412813e-15 pua = -1.50463276905253e-36
+ ub = 7.30246469819168e-19 lub = 9.21800540683538e-25
+ uc = -1.05894772401041e-10 luc = 8.24965543747022e-17
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0145390637694 lu0 = -9.84103748616821e-9
+ a0 = 1.279695175654 la0 = -6.74878816783794e-7
+ keta = 0.00236686763209581 lketa = -4.81460926363185e-08 pketa = 5.04870979341448e-29
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.0789146275940702 lags = 1.01599963925139e-6
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.29522360732579+0*(0.0/sqrt(l*w*mult))} lvoff = 6.12567370176266e-10
+ nfactor = {1.8907185940324+0*(0.1/sqrt(l*w*mult))} lnfactor = -2.71834879839156e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.40966078061423 lpclm = 1.22001243377312e-8
+ pdiblc1 = 0.39
+ pdiblc2 = 0.000215
+ pdiblcb = -0.0485835162604495 lpdiblcb = 9.41769516564709e-8
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 9.98760699558709e-09 lpscbe2 = -1.90232158012223e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -2.1192557782444e-11 lalpha0 = 1.42773752745155e-16 palpha0 = -9.4039548065783e-38
+ alpha1 = -9.78990408614235e-11 lalpha1 = 3.94479678312628e-16 walpha1 = 4.00593428432545e-32 palpha1 = 3.58525777000798e-37
+ beta0 = -0.505055838463804 lbeta0 = 1.39968726718594e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.1264173309365e-10 lagidl = 9.2233955698489e-17
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.431177870254609 lkt1 = -8.66147814024155e-8
+ kt2 = -0.046670102192069 lkt2 = -1.89983007746655e-8
+ at = 65353.85212337 lat = -0.0760016964958941
+ ute = 0.73294808402065 lute = -3.54823748770555e-06 wute = -4.2351647362715e-22 pute = 8.07793566946316e-28
+ ua1 = 4.5307033248294e-09 lua1 = -9.38179145816879e-15
+ ub1 = -2.45594843985464e-18 lub1 = 6.12082028642296e-24
+ uc1 = -2.7031855873761e-10 luc1 = 5.5897494905091e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.40 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.004443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.0461095036822+0*(0.005856/sqrt(l*w*mult))} lvth0 = 4.93666175802686e-8
+ k1 = 0.5454080839698 lk1 = -6.41976508749527e-8
+ k2 = -0.0229531449202714 lk2 = 2.50713315250286e-08 wk2 = 2.64697796016969e-23
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -29678.9552125641 lvsat = 0.108224007437026
+ ua = -2.46780240508459e-10 lua = -1.10389310181221e-15
+ ub = 8.93180803063238e-19 lub = 5.97017342723469e-25
+ uc = -9.8690946200604e-11 luc = 6.81368938639755e-17
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0121160398104 lu0 = -5.01113175378311e-9
+ a0 = 0.823582341107999 la0 = 2.34308228604462e-7
+ keta = -0.0355693011631478 lketa = 2.74735141976547e-8
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.540114866427679 lags = 9.66716775752801e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.28425387944166+0*(0.0/sqrt(l*w*mult))} lvoff = -2.12538080709206e-8
+ nfactor = {1.9294746740774+0*(0.1/sqrt(l*w*mult))} lnfactor = -3.49088846923894e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = -0.32726858 leta0 = 8.1182393672004e-07 peta0 = 4.03896783473158e-28
+ etab = 22.482326763364 letab = -4.49544099258305e-05 wetab = -1.52465930505774e-20 petab = 1.85792520397653e-26
+ dsub = 0.8580014 ldsub = -5.94017514673199e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.20596428508744 lpclm = 4.18236089338114e-7
+ pdiblc1 = 0.40380624592792 lpdiblc1 = -2.75205146454677e-8
+ pdiblc2 = 1.43232999999954e-06 lpdiblc2 = 4.2571255218246e-10
+ pdiblcb = -0.00189449793638372 lpdiblcb = 1.10995724841425e-09 wpdiblcb = -3.30872245021211e-24
+ drout = 0.36191763501608 ldrout = 3.94845105252317e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 1.06879873224826e-08 lpscbe2 = -3.29841630017542e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.19602200021382e-12 lalpha0 = 9.81457458983515e-17
+ alpha1 = 1.0e-10
+ beta0 = 4.1721815058722 lbeta0 = 4.67355773837533e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 2.1743320265992e-10 lagidl = -1.16650862663799e-16
+ bgidl = 802899192.027399 lbgidl = 392.888530362485
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.499503183519999 lkt1 = 4.95806618913891e-8
+ kt2 = -0.0621669880279999 lkt2 = 1.18922306437576e-8
+ at = -10090.728646 lat = 0.0743848532457603
+ ute = -1.6830846545 lute = 1.26773237923172e-6
+ ua1 = -6.0105839752e-10 lua1 = 8.47544189935722e-16 wua1 = -7.88860905221012e-31 pua1 = -7.52316384526264e-37
+ ub1 = 7.16179343459999e-19 lub1 = -2.0230256491387e-25
+ uc1 = -7.3692013666e-11 luc1 = 1.67031784950957e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.41 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.004443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.0191663245768+0*(0.005856/sqrt(l*w*mult))} lvth0 = 2.26029339340689e-8
+ k1 = 0.51047242407276 lk1 = -2.94947323441476e-8
+ k2 = -0.014917698045952 lk2 = 1.70894167977859e-08 wk2 = 6.61744490042422e-24 pk2 = -3.15544362088405e-30
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 69602.3155281761 lvsat = 0.00960414852196073
+ ua = -1.5165106213508e-09 lua = 1.57378335232962e-16
+ ub = 1.5753040065058e-18 lub = -8.05615559377569e-26
+ uc = -5.27318395745652e-11 luc = 2.24839668062795e-17 puc = 4.70197740328915e-38
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.00663341319120002 lu0 = 4.34969606879781e-10
+ a0 = 1.113099680712 la0 = -5.32803464830964e-8
+ keta = -0.00348616462015641 lketa = -4.39588448968729e-9
+ a1 = 0.0
+ a2 = 0.75935673367364 la2 = 4.03725008860941e-8
+ ags = 0.277159512155241 lags = 3.57875223277558e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.272911688847361+0*(0.0/sqrt(l*w*mult))} lvoff = -3.2520436991481e-8
+ nfactor = {1.2567334619324+0*(0.1/sqrt(l*w*mult))} lnfactor = 3.19170563265793e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.49
+ etab = -45.243261151015 letab = 2.2319990121863e-5
+ dsub = 0.231063940416441 ldsub = 2.87432875546143e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.63111242831704 lpclm = -4.07971696129197e-9
+ pdiblc1 = 0.5605837704226 lpdiblc1 = -1.83253587271965e-7
+ pdiblc2 = 0.000274683463070081 lpdiblc2 = 1.54281818160893e-10
+ pdiblcb = 0.220458260914565 lpdiblcb = -2.1976148752307e-07 wpdiblcb = -2.9778502051909e-23 ppdiblcb = 8.67746995743113e-29
+ drout = 0.522027289967841 ldrout = 2.35802100821845e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 5.437709665876e-09 lpscbe2 = 1.91688400668287e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.37476536438882 lbeta0 = 4.98971493524157e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -6.12587401723994e-12 lagidl = 1.05418863444537e-16
+ bgidl = 1394201615.9452 lbgidl = -194.474636807174
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.391504383880001 lkt1 = -5.76986497454084e-8
+ kt2 = -0.0452685267320001 lkt2 = -4.89365310308852e-9
+ at = 55827.0751880002 lat = 0.00890619382090246
+ ute = -0.49488123272 lute = 8.74447686476193e-8
+ ua1 = -4.78189710399998e-11 lua1 = 2.97990444514932e-16
+ ub1 = 6.06412088160001e-19 lub1 = -9.32665790686781e-26
+ uc1 = 1.6366545464e-10 luc1 = -6.87444079011884e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.42 pmos
* DC IV MOS Parameters
+ lmin = 2.5e-07 lmax = 5e-07 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.006443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.951579035816+0*(0.007356/sqrt(l*w*mult))} lvth0 = -1.07404439286061e-8
+ k1 = 0.139138830563601 lk1 = 1.53698240010475e-7
+ k2 = 0.117740448063352 lk2 = -4.83558876874859e-08 wk2 = -1.05879118406788e-22 pk2 = -3.78653234506086e-29
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 70255.1058400003 lvsat = 0.00928210225510606
+ ua = -4.86169000896802e-10 lua = -3.50928339118575e-16
+ ub = 1.0420180418272e-18 lub = 1.82528675304854e-25
+ uc = -7.86051795167599e-12 luc = 3.47238739486536e-19
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.01055413854848 lu0 = -1.49927319943002e-9
+ a0 = 1.49585434488 la0 = -2.42107766994409e-07 wa0 = 3.3881317890172e-21
+ keta = 0.050567389226496 lketa = -3.10625566372871e-08 wketa = -5.29395592033938e-23 pketa = -1.26217744835362e-29
+ a1 = 0.0
+ a2 = 0.88128653265272 la2 = -1.97801022826479e-8
+ ags = 1.097940292214 lags = -4.70471251950699e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.26197424659896+0*(0.0/sqrt(l*w*mult))} lvoff = -3.79162928754222e-8
+ nfactor = {1.1099157291336+0*(0.1/sqrt(l*w*mult))} lnfactor = 3.91601329929288e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.681857840994881 leta0 = -9.46507635607321e-8
+ etab = -0.000870723701341264 letab = 1.99713232889716e-10
+ dsub = 0.0824405601279206 ldsub = 1.02064848739392e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.40264312934008 lpclm = 1.08632870057403e-7
+ pdiblc1 = -0.00365505965855961 lpdiblc1 = 9.51068686826147e-8
+ pdiblc2 = -0.00640266916101695 lpdiblc2 = 3.44847360702275e-09 wpdiblc2 = -3.30872245021211e-24 ppdiblc2 = -1.18329135783152e-30
+ pdiblcb = -0.3225732332316 lpdiblcb = 4.81365837360111e-8
+ drout = 1.40305344137712 ldrout = -1.98841578662105e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 9.4174066817368e-09 lpscbe2 = -4.64517597278732e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 9.8374004106232 lbeta0 = -2.22601954915031e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -2.08500774325672e-09 lagidl = 1.1310102870514e-15 pagidl = 5.64237288394698e-37
+ bgidl = 1000000000.0
+ cgidl = 532.846726441352 lcgidl = -0.000114872138329124
+ egidl = -1.1321491658048 legidl = 6.07866005159808e-07 wegidl = 8.470329472543e-22 pegidl = -1.0097419586829e-28
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.48341565304 lkt1 = -1.23553280405526e-8
+ kt2 = -0.049672987568 lkt2 = -2.72076520317801e-9
+ at = 91080.1031920002 lat = -0.00848546450853488
+ ute = -0.33479019576 lute = 8.46577665584676e-9
+ ua1 = 9.01049146560001e-10 lua1 = -1.70122254885617e-16 wua1 = 1.57772181044202e-30
+ ub1 = 4.4136286032e-19 lub1 = -1.18415231045482e-26
+ uc1 = 4.74074714316e-11 luc1 = -1.13899269811227e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.24e-6
+ sbref = 1.24e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.43 pmos
* DC IV MOS Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.006443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.785792300714288+0*(0.007356/sqrt(l*w*mult))} lvth0 = -5.10826564747865e-8
+ k1 = 0.109830032788 lk1 = 1.60830184243594e-7
+ k2 = 0.140327289931343 lk2 = -5.38521246139592e-8
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 199357.877371429 lvsat = -0.0221335079638087
+ ua = -1.20274672320286e-09 lua = -1.76557749328064e-16
+ ub = 1.15786067182572e-18 lub = 1.54339761406273e-25
+ uc = -2.29894954758249e-11 luc = 4.02869387225787e-18
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.00679047121600002 lu0 = -5.83429918079004e-10
+ a0 = -0.464755997999996 la0 = 2.34983232621324e-7
+ keta = -0.327136074690686 lketa = 6.08470488653921e-8
+ a1 = 0.0
+ a2 = 1.117265914878 la2 = -7.72028531945829e-8
+ ags = 0.04929956616715 lags = 2.0812701179972e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.218487508549716+0*(0.0/sqrt(l*w*mult))} lvoff = -4.84982687388494e-8
+ nfactor = {1.36988594933716+0*(0.1/sqrt(l*w*mult))} lnfactor = 3.28340696485398e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.567449993717428 leta0 = -6.68109868199315e-8
+ etab = 0.193850720008982 letab = -4.71834134366929e-08 wetab = 4.01182597088218e-23 petab = 8.97329279688901e-30
+ dsub = 1.07184049999343 ldsub = -1.38693753827601e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.38934427018857 lpclm = -1.31469012154386e-7
+ pdiblc1 = 0.898253486238859 lpdiblc1 = -1.24361753058971e-7
+ pdiblc2 = 0.0170353361227257 lpdiblc2 = -2.25488372271263e-9
+ pdiblcb = -0.433203011048126 lpdiblcb = 7.50570126103288e-8
+ drout = -0.439476576346854 ldrout = 2.49515990790812e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 8.60635267050003e-09 lpscbe2 = 1.50908501258468e-16
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 9.76940471184574 lbeta0 = -2.06056017565909e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 8.16250109563772e-09 lagidl = -1.36259801878749e-15
+ bgidl = 1000000000.0
+ cgidl = -531.595451576256 lcgidl = 0.000144147092385325
+ egidl = 4.50053273501714 legidl = -7.62779543222403e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.376180031714286 lkt1 = -3.84498296627094e-8
+ kt2 = 0.0904601689714282 lkt2 = -3.68204872491695e-8
+ at = 26226.478514286 lat = 0.00729588681329074
+ ute = -0.3
+ ua1 = 3.68606868285714e-10 lua1 = -4.05588157749091e-17
+ ub1 = 3.927e-19
+ uc1 = 6.0045e-13
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.44 pmos
* DC IV MOS Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.006443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-3.26380050227181+0*(0.007356/sqrt(l*w*mult))} lvth0 = 3.78450329166792e-07 wvth0 = 4.32374301974468e-06 pvth0 = -7.49468967556504e-13
+ k1 = -4.6307136029321 lk1 = 9.82546536972046e-07 wk1 = 7.42601738700357e-06 pk1 = -1.28721100182843e-12
+ k2 = 1.02422191607785 lk2 = -2.07064651320942e-07 wk2 = -1.15912305740656e-06 pk2 = 2.00920072524738e-13
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 363519.32933208 lvsat = -0.0505889257237641 wvsat = -0.271997448857645 pvsat = 4.71474937900866e-8
+ ua = 1.03960618389328e-08 lua = -2.18707202787153e-15 wua = -1.93579282067587e-14 pua = 3.35546455950314e-21
+ ub = -3.57142310780033e-18 lub = 9.74104353199095e-25 wub = 6.72394316230623e-24 pub = -1.16551485986784e-30
+ uc = 6.41418596172956e-13 luc = -6.74415111540877e-20 wuc = 6.55503634637616e-19 puc = -1.13623689020815e-25
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.046625333803371 lu0 = -7.48832532924873e-09 wu0 = -6.94985774249307e-08 pu0 = 1.20467444136826e-14
+ a0 = 8.58968829925363 la0 = -1.33449603297603e-06 wa0 = -1.26394969896403e-05 pa0 = 2.19090512919027e-12
+ keta = 2.04794846789243 lketa = -3.5084535557688e-07 wketa = -3.5336991662667e-06 pketa = 6.12524346082338e-13
+ a1 = 0.0
+ a2 = -0.893484834715334 la2 = 2.71336660238426e-7
+ ags = 37.545363627095 lags = -6.29136574039339e-06 wags = -6.27816221301311e-05 pags = 1.08824408167927e-11
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-3.92087664490584+0*(0.0/sqrt(l*w*mult))} lvoff = 5.93266459378849e-07 wvoff = 5.79962510539864e-06 pvoff = -1.00529541651959e-12
+ nfactor = {41.9938193494667+0*(0.1/sqrt(l*w*mult))} lnfactor = -6.71333067122626e-06 wnfactor = -7.78511966309952e-05 pnfactor = 1.34945707216235e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.225074950427021 leta0 = -7.46438156605941e-09 weta0 = -1.05802190212116e-06 peta0 = 1.83395400469877e-13
+ etab = -1.36540444630799 letab = 2.23094758582359e-07 wetab = 1.87075980821804e-06 petab = -3.24273763636898e-13
+ dsub = 0.318486163890462 ldsub = -8.10881991618481e-09 wdsub = 1.58254023669715e-08 pdsub = -2.7431435954861e-15
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.354485082557115 lpclm = 1.70802880191845e-07 wpclm = 2.95157094618367e-06 ppclm = -5.11619404669587e-13
+ pdiblc1 = 0.95148729129 lpdiblc1 = -1.33589194358926e-7
+ pdiblc2 = 0.0212117343376134 lpdiblc2 = -2.97881223648482e-9
+ pdiblcb = 0.763376357191859 lpdiblcb = -1.32355661921654e-07 wpdiblcb = -1.3221774355697e-06 ppdiblcb = 2.29183592326781e-13
+ drout = 1.0
+ pscbe1 = 1369148945.55987 lpscbe1 = -98.6551399254558 wpscbe1 = -984.4809492204 ppscbe1 = 0.000170647958775967
+ pscbe2 = 1.09522527291816e-08 lpscbe2 = -2.55725123113284e-16 wpscbe2 = -1.27679985792491e-15 ppscbe2 = 2.21317933772982e-22
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 16.3849219927818 lbeta0 = -1.35277655200882e-06 wbeta0 = -4.87962787989939e-06 pbeta0 = 8.45824937445994e-13
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 4.50812115916652e-09 lagidl = -7.29155109359447e-16 wagidl = -7.11547126116867e-15 pagidl = 1.23338155746846e-21
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.0640181706666674 lkt1 = -9.25593423329808e-8
+ kt2 = -0.131324749333333 lkt2 = 1.62326691994133e-9
+ at = 615462.065218183 lat = -0.0948410313147893 wat = -0.705986371733274 pat = 1.22374265703502e-7
+ ute = -0.718403621999999 lute = 7.25252470302358e-8
+ ua1 = 8.98188337989136e-10 lua1 = -1.32355408570361e-16 wua1 = -1.56962326948797e-15 pua1 = 2.72075358286506e-22
+ ub1 = 5.46403897747175e-20 lub1 = 5.85985767172297e-26 wub1 = 7.81370639380857e-25 pub1 = -1.35441223888999e-31
+ uc1 = -2.73406652366667e-11 luc1 = 4.84325703289333e-18 wuc1 = 1.23259516440783e-32 puc1 = -2.93873587705572e-39
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.45 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 1.65e-06 wmax = 1.68e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.004443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.034517+0*(0.005856/sqrt(l*w*mult))}
+ k1 = 0.42302944
+ k2 = 0.023080264
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 53438.0
+ ua = -1.9280657e-10
+ ub = 9.7328962e-19
+ uc = -9.8608028e-11
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0126711
+ a0 = 1.118778
+ keta = 4.9707517e-6
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.17518243
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.29720858+0*(0.0/sqrt(l*w*mult))}
+ nfactor = {1.911951+0*(0.1/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.14877095
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00019189
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 757128280.0
+ pscbe2 = 9.873241e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.7815831e-11
+ alpha1 = 6.3056523e-17
+ beta0 = 9.6797043
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 1352540500.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.4443203
+ kt2 = -0.052664618
+ at = 90000.0
+ ute = -0.17124159
+ ua1 = 2.1098632e-9
+ ub1 = -7.3847396e-19
+ uc1 = 1.1059776e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.46 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 1.65e-06 wmax = 1.68e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.004443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.034517+0*(0.005856/sqrt(l*w*mult))}
+ k1 = 0.42302944
+ k2 = 0.023080264
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 53438.0
+ ua = -1.9280657e-10
+ ub = 9.7328962e-19
+ uc = -9.8608028e-11
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0126711
+ a0 = 1.118778
+ keta = 4.9707517e-6
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.17518243
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.29720858+0*(0.0/sqrt(l*w*mult))}
+ nfactor = {1.911951+0*(0.1/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.14877095
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00019189
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 757128280.0
+ pscbe2 = 9.873241e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.7815831e-11
+ alpha1 = 6.3056523e-17
+ beta0 = 9.6797043
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 1352540500.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.4443203
+ kt2 = -0.052664618
+ at = 90000.0
+ ute = -0.17124159
+ ua1 = 2.1098632e-9
+ ub1 = -7.3847396e-19
+ uc1 = 1.1059776e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.47 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 1.65e-06 wmax = 1.68e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.004443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.03968537770652+0*(0.005856/sqrt(l*w*mult))} lvth0 = 4.13125899196556e-8
+ k1 = 0.390669914700908 lk1 = 2.5866062323523e-7
+ k2 = 0.0351772658317135 lk2 = -9.66954244275032e-8
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 77014.5327768419 lvsat = -0.188455195353377
+ ua = -9.89907109822339e-11 lua = -7.49901870889346e-16
+ ub = 9.85477846643298e-19 lub = -9.74246151805995e-26
+ uc = -1.11957558265435e-10 luc = 1.06707307552853e-16
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0132665066958 lu0 = -4.75928696699256e-9
+ a0 = 1.126848536098 la0 = -6.45105228724895e-8
+ keta = 0.00968353076963805 lketa = -7.73640015766657e-08 wketa = 7.65142066611551e-24 pketa = -8.36192559534273e-29
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.0172899885681765 lags = 1.26208765200977e-6
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.299343388544763+0*(0.0/sqrt(l*w*mult))} lvoff = 1.70642462635792e-8
+ nfactor = {2.00110676335524+0*(0.1/sqrt(l*w*mult))} lnfactor = -7.12652151146605e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.114734399685773 lpclm = 2.1062873248466e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 0.000168818489704996 lpdiblc2 = 1.84418379958404e-10
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 714327962.849655 lpscbe1 = 342.117401489872
+ pscbe2 = 1.02346458760092e-08 lpscbe2 = -2.88883132878909e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.10658131246379e-11 lalpha0 = -2.59782056161903e-17
+ alpha1 = -8.83803561262885e-13 lalpha1 = 7.06504462287933e-18 walpha1 = 1.85521220424177e-33 palpha1 = -4.32200803793546e-39
+ beta0 = 16.3482835524883 lbeta0 = -5.33042079449266e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 6.43208327881965e-11 lagidl = 2.85195643082482e-16
+ bgidl = 1704493843.79724 lbgidl = -2813.28203720157
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.435787145678042 lkt1 = -6.82083867015442e-8
+ kt2 = -0.0538995747481872 lkt2 = 9.87142670363705e-9
+ at = 133605.523841314 lat = -0.348553690730682
+ ute = -0.186865964192179 lute = 1.24890903956579e-7
+ ua1 = 2.03850284894073e-09 lua1 = 5.70407405815369e-16
+ ub1 = -5.540650054973e-19 lub1 = -1.47404310356667e-24
+ uc1 = 3.51135925346025e-10 luc1 = -1.92270285751065e-15
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.48 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 1.65e-06 wmax = 1.68e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.004443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.0373096643247+0*(0.005856/sqrt(l*w*mult))} lvth0 = 3.18255633950442e-8
+ k1 = 0.397876315328929 lk1 = 2.29883029764097e-7
+ k2 = 0.0322306662092167 lk2 = -8.4928656184203e-08 pk2 = -8.07793566946316e-28
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 35013.0233625527 lvsat = -0.0207289717519412
+ ua = 2.2530214708256e-10 lua = -2.04491286412813e-15
+ ub = 7.30246469819167e-19 lub = 9.21800540683505e-25
+ uc = -1.05894772401042e-10 luc = 8.24965543747053e-17
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0145390637694001 lu0 = -9.8410374861681e-9
+ a0 = 1.279695175654 la0 = -6.74878816783818e-7
+ keta = 0.00236686763209581 lketa = -4.8146092636319e-8
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.0789146275940666 lags = 1.0159996392514e-6
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.295223607325795+0*(0.0/sqrt(l*w*mult))} lvoff = 6.12567370160172e-10
+ nfactor = {1.89071859403239+0*(0.1/sqrt(l*w*mult))} lnfactor = -2.71834879839183e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.409660780614232 lpclm = 1.22001243377414e-8
+ pdiblc1 = 0.39
+ pdiblc2 = 0.000215
+ pdiblcb = -0.0485835162604493 lpdiblcb = 9.41769516564715e-8
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 9.98760699558733e-09 lpscbe2 = -1.90232158012228e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -2.11925577824438e-11 lalpha0 = 1.42773752745155e-16 palpha0 = -1.50463276905253e-36
+ alpha1 = -9.78990408614231e-11 lalpha1 = 3.94479678312631e-16 walpha1 = 2.46519032881566e-31 palpha1 = -2.82118644197349e-37
+ beta0 = -0.505055838463818 lbeta0 = 1.39968726718595e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.12641733093649e-10 lagidl = 9.22339556984973e-17
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.431177870254608 lkt1 = -8.66147814024206e-8
+ kt2 = -0.0466701021920688 lkt2 = -1.89983007746662e-8
+ at = 65353.8521233695 lat = -0.0760016964958936
+ ute = 0.732948084020652 lute = -3.54823748770557e-06 wute = -6.7762635780344e-21 pute = 1.29246970711411e-26
+ ua1 = 4.53070332482936e-09 lua1 = -9.38179145816882e-15 wua1 = 5.04870979341448e-29
+ ub1 = -2.45594843985465e-18 lub1 = 6.12082028642299e-24 wub1 = 2.35098870164458e-38
+ uc1 = -2.7031855873761e-10 luc1 = 5.58974949050908e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.49 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 1.65e-06 wmax = 1.68e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.004443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.04610950368219+0*(0.005856/sqrt(l*w*mult))} lvth0 = 4.93666175802737e-8
+ k1 = 0.545408083969797 lk1 = -6.41976508749536e-8
+ k2 = -0.0229531449202711 lk2 = 2.50713315250286e-8
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -29678.9552125637 lvsat = 0.108224007437025 pvsat = -8.470329472543e-22
+ ua = -2.46780240508439e-10 lua = -1.1038931018122e-15
+ ub = 8.93180803063207e-19 lub = 5.97017342723471e-25
+ uc = -9.86909462006028e-11 luc = 6.81368938639742e-17 wuc = 1.57772181044202e-30
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0121160398103999 lu0 = -5.01113175378287e-9
+ a0 = 0.823582341107993 la0 = 2.34308228604449e-7
+ keta = -0.0355693011631475 lketa = 2.74735141976551e-8
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.540114866427672 lags = 9.66716775752742e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.284253879441657+0*(0.0/sqrt(l*w*mult))} lvoff = -2.12538080709266e-8
+ nfactor = {1.92947467407737+0*(0.1/sqrt(l*w*mult))} lnfactor = -3.49088846923897e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = -0.327268580000002 leta0 = 8.11823936720047e-7
+ etab = 22.482326763364 letab = -4.49544099258304e-05 wetab = 1.01643953670516e-19 petab = 2.81112161297318e-25
+ dsub = 0.858001399999992 ldsub = -5.94017514673198e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.205964285087447 lpclm = 4.18236089338124e-7
+ pdiblc1 = 0.40380624592791 lpdiblc1 = -2.75205146454694e-8
+ pdiblc2 = 1.43232999999868e-06 lpdiblc2 = 4.2571255218246e-10
+ pdiblcb = -0.00189449793638372 lpdiblcb = 1.10995724841424e-9
+ drout = 0.36191763501607 ldrout = 3.94845105252322e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 1.06879873224827e-08 lpscbe2 = -3.29841630017526e-15 wpscbe2 = 2.01948391736579e-28
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.19602200021331e-12 lalpha0 = 9.81457458983526e-17
+ alpha1 = 1.0e-10
+ beta0 = 4.17218150587212 lbeta0 = 4.6735577383753e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 2.17433202659919e-10 lagidl = -1.16650862663801e-16
+ bgidl = 802899192.027405 lbgidl = 392.888530362499
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.499503183519998 lkt1 = 4.95806618913848e-8
+ kt2 = -0.0621669880280002 lkt2 = 1.18922306437576e-8
+ at = -10090.7286460004 lat = 0.0743848532457601
+ ute = -1.68308465449999 lute = 1.26773237923172e-6
+ ua1 = -6.01058397519999e-10 lua1 = 8.47544189935723e-16 wua1 = -6.31088724176809e-30 pua1 = 6.01853107621011e-36
+ ub1 = 7.16179343459997e-19 lub1 = -2.02302564913869e-25
+ uc1 = -7.36920136659996e-11 luc1 = 1.67031784950959e-16 wuc1 = -3.94430452610506e-31 puc1 = -7.52316384526264e-37
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.50 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 1.65e-06 wmax = 1.68e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.004443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.0191663245768+0*(0.005856/sqrt(l*w*mult))} lvth0 = 2.26029339340765e-8
+ k1 = 0.510472424072759 lk1 = -2.94947323441447e-8
+ k2 = -0.0149176980459521 lk2 = 1.7089416797786e-08 pk2 = -5.04870979341448e-29
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 69602.3155281767 lvsat = 0.00960414852196134
+ ua = -1.51651062135081e-09 lua = 1.57378335232956e-16
+ ub = 1.57530400650579e-18 lub = -8.05615559377525e-26
+ uc = -5.27318395745649e-11 luc = 2.24839668062795e-17
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.00663341319120003 lu0 = 4.3496960687982e-10
+ a0 = 1.11309968071201 la0 = -5.32803464831032e-8
+ keta = -0.00348616462015638 lketa = -4.39588448968723e-9
+ a1 = 0.0
+ a2 = 0.759356733673641 la2 = 4.03725008861001e-8
+ ags = 0.277159512155237 lags = 3.57875223277557e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.272911688847365+0*(0.0/sqrt(l*w*mult))} lvoff = -3.25204369914785e-8
+ nfactor = {1.25673346193241+0*(0.1/sqrt(l*w*mult))} lnfactor = 3.1917056326579e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.49
+ etab = -45.2432611510153 letab = 2.2319990121863e-5
+ dsub = 0.231063940416441 ldsub = 2.87432875546154e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.631112428317024 lpclm = -4.07971696129197e-9
+ pdiblc1 = 0.560583770422603 lpdiblc1 = -1.83253587271961e-7
+ pdiblc2 = 0.00027468346307008 lpdiblc2 = 1.54281818160896e-10
+ pdiblcb = 0.220458260914567 lpdiblcb = -2.1976148752307e-07 wpdiblcb = 5.82335151237331e-22 ppdiblcb = -2.39813715187188e-28
+ drout = 0.522027289967838 ldrout = 2.35802100821851e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 5.43770966587597e-09 lpscbe2 = 1.91688400668291e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.37476536438874 lbeta0 = 4.98971493524225e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -6.12587401724014e-12 lagidl = 1.05418863444536e-16
+ bgidl = 1394201615.94521 lbgidl = -194.474636807165
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.391504383879997 lkt1 = -5.76986497454101e-8
+ kt2 = -0.0452685267320003 lkt2 = -4.89365310308889e-9
+ at = 55827.0751879988 lat = 0.00890619382090296
+ ute = -0.494881232719997 lute = 8.74447686476193e-8
+ ua1 = -4.78189710399998e-11 lua1 = 2.97990444514927e-16 pua1 = 3.00926553810506e-36
+ ub1 = 6.06412088159995e-19 lub1 = -9.32665790686762e-26
+ uc1 = 1.63665454639999e-10 luc1 = -6.87444079011878e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.51 pmos
* DC IV MOS Parameters
+ lmin = 2.5e-07 lmax = 5e-07 wmin = 1.65e-06 wmax = 1.68e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.006443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.951579035815996+0*(0.007356/sqrt(l*w*mult))} lvth0 = -1.07404439286048e-8
+ k1 = 0.13913883056361 lk1 = 1.53698240010471e-7
+ k2 = 0.117740448063352 lk2 = -4.83558876874858e-08 wk2 = 4.2351647362715e-22 pk2 = -2.01948391736579e-28
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 70255.1058399994 lvsat = 0.00928210225510595
+ ua = -4.86169000896822e-10 lua = -3.50928339118571e-16
+ ub = 1.04201804182721e-18 lub = 1.82528675304856e-25
+ uc = -7.86051795167597e-12 luc = 3.47238739486555e-19
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0105541385484801 lu0 = -1.49927319943001e-9
+ a0 = 1.49585434488003 la0 = -2.4210776699441e-7
+ keta = 0.0505673892264957 lketa = -3.1062556637287e-08 wketa = -4.2351647362715e-22 pketa = -2.01948391736579e-28
+ a1 = 0.0
+ a2 = 0.881286532652723 la2 = -1.9780102282645e-8
+ ags = 1.09794029221402 lags = -4.70471251950711e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.26197424659896+0*(0.0/sqrt(l*w*mult))} lvoff = -3.79162928754216e-8
+ nfactor = {1.10991572913366+0*(0.1/sqrt(l*w*mult))} lnfactor = 3.91601329929288e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.68185784099488 leta0 = -9.46507635607311e-8
+ etab = -0.000870723701341267 letab = 1.99713232889717e-10
+ dsub = 0.082440560127921 ldsub = 1.02064848739392e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.402643129340092 lpclm = 1.08632870057402e-7
+ pdiblc1 = -0.00365505965856272 lpdiblc1 = 9.51068686826138e-8
+ pdiblc2 = -0.00640266916101692 lpdiblc2 = 3.44847360702274e-09 wpdiblc2 = 5.29395592033938e-23 ppdiblc2 = 2.52435489670724e-29
+ pdiblcb = -0.322573233231598 lpdiblcb = 4.81365837360113e-8
+ drout = 1.40305344137712 ldrout = -1.98841578662106e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 9.4174066817369e-09 lpscbe2 = -4.64517597278543e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 9.83740041062333 lbeta0 = -2.22601954914976e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -2.0850077432567e-09 lagidl = 1.1310102870514e-15 wagidl = -6.31088724176809e-30 pagidl = 9.02779661431517e-36
+ bgidl = 1000000000.0
+ cgidl = 532.846726441356 lcgidl = -0.000114872138329124
+ egidl = -1.1321491658048 legidl = 6.07866005159807e-07 pegidl = 3.23117426778526e-27
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.483415653040005 lkt1 = -1.23553280405532e-8
+ kt2 = -0.049672987568 lkt2 = -2.72076520317804e-9
+ at = 91080.1031920016 lat = -0.0084854645085346
+ ute = -0.334790195760007 lute = 8.46577665584697e-9
+ ua1 = 9.01049146560002e-10 lua1 = -1.70122254885617e-16 pua1 = -3.00926553810506e-36
+ ub1 = 4.41362860320004e-19 lub1 = -1.18415231045478e-26
+ uc1 = 4.74074714316003e-11 luc1 = -1.13899269811226e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.24e-6
+ sbref = 1.24e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.52 pmos
* DC IV MOS Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 1.65e-06 wmax = 1.68e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.006443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.785792300714292+0*(0.007356/sqrt(l*w*mult))} lvth0 = -5.10826564747874e-8
+ k1 = 0.109830032788011 lk1 = 1.608301842436e-7
+ k2 = 0.140327289931342 lk2 = -5.38521246139583e-8
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 199357.87737143 lvsat = -0.0221335079638085
+ ua = -1.20274672320286e-09 lua = -1.76557749328069e-16
+ ub = 1.15786067182574e-18 lub = 1.54339761406275e-25
+ uc = -2.29894954758248e-11 luc = 4.02869387225789e-18
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.00679047121599996 lu0 = -5.83429918079021e-10
+ a0 = -0.464755998000015 la0 = 2.34983232621319e-7
+ keta = -0.327136074690687 lketa = 6.08470488653919e-08 wketa = -3.3881317890172e-21
+ a1 = 0.0
+ a2 = 1.11726591487798 la2 = -7.72028531945821e-8
+ ags = 0.04929956616715 lags = 2.08127011799721e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.218487508549714+0*(0.0/sqrt(l*w*mult))} lvoff = -4.84982687388487e-8
+ nfactor = {1.36988594933712+0*(0.1/sqrt(l*w*mult))} lnfactor = 3.28340696485388e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.567449993717432 leta0 = -6.6810986819931e-8
+ etab = 0.193850720008983 letab = -4.71834134366926e-08 wetab = -7.17992771696028e-22 petab = 1.73549399148623e-29
+ dsub = 1.07184049999343 ldsub = -1.386937538276e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.38934427018856 lpclm = -1.31469012154386e-7
+ pdiblc1 = 0.898253486238843 lpdiblc1 = -1.24361753058972e-7
+ pdiblc2 = 0.0170353361227258 lpdiblc2 = -2.25488372271259e-9
+ pdiblcb = -0.433203011048128 lpdiblcb = 7.50570126103286e-8
+ drout = -0.439476576346863 ldrout = 2.49515990790809e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 8.60635267050024e-09 lpscbe2 = 1.50908501258494e-16
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 9.76940471184571 lbeta0 = -2.06056017565902e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 8.16250109563776e-09 lagidl = -1.36259801878749e-15
+ bgidl = 1000000000.0
+ cgidl = -531.595451576264 lcgidl = 0.000144147092385324
+ egidl = 4.50053273501715 legidl = -7.62779543222397e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.376180031714298 lkt1 = -3.84498296627107e-8
+ kt2 = 0.0904601689714273 lkt2 = -3.68204872491697e-8
+ at = 26226.4785142858 lat = 0.00729588681329041
+ ute = -0.3
+ ua1 = 3.68606868285714e-10 lua1 = -4.05588157749085e-17
+ ub1 = 3.927e-19
+ uc1 = 6.0045e-13
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.53 pmos
* DC IV MOS Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 1.65e-06 wmax = 1.68e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.006443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {4.01114330042014+0*(0.007356/sqrt(l*w*mult))} lvth0 = -8.82573879704224e-07 wvth0 = -8.26003427840006e-06 pvth0 = 1.43177782174931e-12
+ k1 = -0.337578251893376 lk1 = 2.38383041493692e-7
+ k2 = -0.874877798950216 lk2 = 1.22121495082591e-07 wk2 = 2.12582986168546e-06 pk2 = -3.68487096564832e-13
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 4323.3989690505 lvsat = 0.0116733784535028 wvsat = 0.34931890995955 pvsat = -6.0550241214568e-8
+ ua = 1.74652235615312e-09 lua = -6.87778153005483e-16 wua = -4.39645475282877e-15 pua = 7.62072673945822e-22
+ ub = 3.02291348007139e-18 lub = -1.68944762269392e-25 wub = -4.68255911473907e-24 pub = 8.11665431830666e-31
+ uc = 1.02037890288087e-12 luc = -1.33129732798224e-19
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0113547034459058 lu0 = -1.37458480434643e-09 wu0 = -8.48947967502222e-09 pu0 = 1.47154942790896e-15
+ a0 = 1.28253178214936 la0 = -6.78881366141971e-8
+ keta = 0.00504336546346629 lketa = 3.26772906795149e-9
+ a1 = 0.0
+ a2 = -0.893484834715338 la2 = 2.71336660238429e-7
+ ags = 1.25
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-2.73636761547218+0*(0.0/sqrt(l*w*mult))} lvoff = 3.87946033234868e-07 wvoff = 3.75072985090612e-06 pvoff = -6.50144010896371e-13
+ nfactor = {49.0978064798815+0*(0.1/sqrt(l*w*mult))} lnfactor = -7.94472159243803e-06 wnfactor = -9.01392629587307e-05 pnfactor = 1.56245595627403e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = -0.386589552018002 leta0 = 9.85603199587557e-8
+ etab = -0.283879229302801 letab = 3.56253405171125e-8
+ dsub = 0.327635158675349 ldsub = -9.69468837420422e-9
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.35187956888265 lpclm = -1.24974955759423e-7
+ pdiblc1 = 0.951487291290007 lpdiblc1 = -1.33589194358926e-7
+ pdiblc2 = 0.0212117343376135 lpdiblc2 = -2.97881223648482e-9
+ pdiblcb = -0.00100196205692768 lpdiblcb = 1.40147180292528e-10
+ drout = 1.0
+ pscbe1 = 800000000.0
+ pscbe2 = 1.02141081328798e-08 lpscbe2 = -1.27776615079535e-16
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 13.5639074624669 lbeta0 = -8.63787535353047e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 3.94518992804005e-10 lagidl = -1.61115370464976e-17
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.0640181706666567 lkt1 = -9.25593423329778e-8
+ kt2 = -0.131324749333331 lkt2 = 1.62326691994176e-9
+ at = 207316.636533339 lat = -0.0240939189974152
+ ute = -0.718403622000011 lute = 7.25252470302352e-8
+ ua1 = -9.24357266666552e-12 lua1 = 2.4937023958895e-17
+ ub1 = 5.0636703399999e-19 lub1 = -1.97028163394924e-26
+ uc1 = -2.73406652366669e-11 luc1 = 4.84325703289333e-18 puc1 = 1.17549435082229e-38
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.54 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 1.26e-06 wmax = 1.65e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.004443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.13241955778733+0*(0.005856/sqrt(l*w*mult))} wvth0 = 1.66409108959069e-7
+ k1 = 0.192177033644933 wk1 = 3.92389577053255e-7
+ k2 = 0.10889696070478 wk2 = -1.45866260853715e-7
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 47393.65057134 wvsat = 0.0102738357954393
+ ua = 3.84222479981006e-09 wua = -6.85851309758997e-15
+ ub = -1.01712351918573e-18 wub = 3.38318920810846e-24
+ uc = -2.9907055997136e-10 wuc = 3.40734625110569e-16
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0309163958791707 wu0 = -3.10122993573125e-8
+ a0 = 0.68344991754 wa0 = 7.3994551260234e-7
+ keta = -0.0222783333676765 wketa = 3.78758723671381e-8
+ a1 = 0.0
+ a2 = 0.8
+ ags = -0.0822918634785329 wags = 4.37639922040647e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.289281852289933+0*(0.0/sqrt(l*w*mult))} wvoff = -1.347339359671e-8
+ nfactor = {2.381769632056+0*(0.1/sqrt(l*w*mult))} wnfactor = -7.98570555251856e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.642546162609021 wpclm = -8.39290566185525e-7
+ pdiblc1 = 0.39
+ pdiblc2 = -0.00107066232286653 wpdiblc2 = 2.14601346288427e-9
+ pdiblcb = 0.646662666666666 wpdiblcb = -1.14165337869787e-6
+ drout = 0.56
+ pscbe1 = 613201011.8902 wpscbe1 = 244.639251336941
+ pscbe2 = 6.85502405793333e-09 wpscbe2 = 5.13019070518567e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 7.76469737917133e-11 walpha0 = -1.01697518277301e-16
+ alpha1 = 2.7482008494454e-16 walpha1 = -3.59943462659449e-22
+ beta0 = -58.562215686586 wbeta0 = 0.000115993671210224
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -5.68598976745332e-11 wagidl = 2.66621387565086e-16
+ bgidl = 2536481961.69 wbgidl = -2012.39526476418
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.104157749960667 wkt1 = -5.78188641161467e-7
+ kt2 = -0.05327118983764 wkt2 = 1.03101574976824e-9
+ at = 358665.066666667 wat = -0.456661351479146
+ ute = 3.48347113841513 wute = -6.21206945336434e-6
+ ua1 = 1.00553410450693e-08 wua1 = -1.35052639924294e-14
+ ub1 = -4.87864951938746e-18 wub1 = 7.03723111369948e-24
+ uc1 = 4.544979784468e-10 wuc1 = -5.84541713883244e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.55 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 1.26e-06 wmax = 1.65e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.004443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.13241955778733+0*(0.005856/sqrt(l*w*mult))} wvth0 = 1.66409108959069e-7
+ k1 = 0.192177033644934 wk1 = 3.92389577053254e-7
+ k2 = 0.10889696070478 wk2 = -1.45866260853715e-7
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 47393.65057134 wvsat = 0.0102738357954394
+ ua = 3.84222479981006e-09 wua = -6.85851309758997e-15
+ ub = -1.01712351918573e-18 wub = 3.38318920810846e-24
+ uc = -2.9907055997136e-10 wuc = 3.4073462511057e-16
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0309163958791707 wu0 = -3.10122993573125e-8
+ a0 = 0.683449917539999 wa0 = 7.39945512602341e-7
+ keta = -0.0222783333676765 wketa = 3.78758723671381e-8
+ a1 = 0.0
+ a2 = 0.8
+ ags = -0.0822918634785332 wags = 4.37639922040648e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.289281852289933+0*(0.0/sqrt(l*w*mult))} wvoff = -1.347339359671e-8
+ nfactor = {2.381769632056+0*(0.1/sqrt(l*w*mult))} wnfactor = -7.98570555251856e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.642546162609021 wpclm = -8.39290566185525e-7
+ pdiblc1 = 0.39
+ pdiblc2 = -0.00107066232286653 wpdiblc2 = 2.14601346288427e-9
+ pdiblcb = 0.646662666666666 wpdiblcb = -1.14165337869787e-6
+ drout = 0.56
+ pscbe1 = 613201011.8902 wpscbe1 = 244.639251336941
+ pscbe2 = 6.85502405793333e-09 wpscbe2 = 5.13019070518566e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 7.76469737917133e-11 walpha0 = -1.01697518277301e-16
+ alpha1 = 2.7482008494454e-16 walpha1 = -3.59943462659448e-22
+ beta0 = -58.562215686586 wbeta0 = 0.000115993671210224
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -5.68598976745332e-11 wagidl = 2.66621387565086e-16
+ bgidl = 2536481961.69 wbgidl = -2012.39526476418
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.104157749960666 wkt1 = -5.78188641161466e-7
+ kt2 = -0.05327118983764 wkt2 = 1.03101574976829e-9
+ at = 358665.066666667 wat = -0.456661351479146
+ ute = 3.48347113841513 wute = -6.21206945336434e-6
+ ua1 = 1.00553410450693e-08 wua1 = -1.35052639924294e-14
+ ub1 = -4.87864951938746e-18 wub1 = 7.03723111369948e-24
+ uc1 = 4.544979784468e-10 wuc1 = -5.84541713883244e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.56 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 1.26e-06 wmax = 1.65e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.004443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.14806250351302+0*(0.005856/sqrt(l*w*mult))} lvth0 = 1.25039352501092e-07 wvth0 = 1.84213174248057e-07 pvth0 = -1.42313911628938e-13
+ k1 = -0.089708682303987 lk1 = 2.25320780495171e-06 wk1 = 8.16519773306009e-07 pk1 = -3.3902160146546e-12
+ k2 = 0.204376147370209 lk2 = -7.63197410981866e-07 wk2 = -2.87594479143781e-07 pk2 = 1.13288155293028e-12
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 108265.231128122 lvsat = -0.486567117984583 wvsat = -0.0531181307671393 pvsat = 5.06713415219389e-7
+ ua = 6.15438713277867e-09 lua = -1.84818950382866e-14 wua = -1.06291302135854e-14 pua = 3.01398170767368e-20
+ ub = -1.92887118191961e-18 lub = 7.28790723894186e-24 wub = 4.95364202937741e-24 pub = -1.25531602134563e-29
+ uc = -4.09735559396951e-10 luc = 8.84582745178557e-16 wuc = 5.06145834754887e-16 puc = -1.32218770767589e-21
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0421160363720325 lu0 = -8.95225119379315e-08 wu0 = -4.90367630408447e-08 pu0 = 1.44075630491199e-13
+ a0 = 0.471748982998644 la0 = 1.69219712470496e-06 wa0 = 1.11350035560412e-06 pa0 = -2.98595012165015e-12
+ keta = 0.00844478630403462 lketa = -2.45580279950436e-07 wketa = 2.10554624320277e-09 pketa = 2.85924307078845e-13
+ a1 = 0.0
+ a2 = 0.8
+ ags = -0.595762931923631 lags = 4.1043478033028e-06 wags = 1.04203191979317e-06 pags = -4.83110952253113e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.235768414400914+0*(0.0/sqrt(l*w*mult))} lvoff = -4.27750996588934e-07 wvoff = -1.08061066416212e-07 pvoff = 7.56071239479694e-13
+ nfactor = {3.81134522329346+0*(0.1/sqrt(l*w*mult))} lnfactor = -1.14270808973109e-05 wnfactor = -3.07693870241999e-06 pnfactor = 1.82117666887487e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.384311688958626 lpclm = 8.20802188553403e-06 wpclm = 4.58211894738672e-07 ppclm = -1.03713757259989e-11
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00040472403201286 lpdiblc2 = -1.17932618151389e-08 wpdiblc2 = -4.00978605474555e-10 ppdiblc2 = 2.03589684857112e-14
+ pdiblcb = 0.646662666666666 wpdiblcb = -1.14165337869787e-6
+ drout = 0.56
+ pscbe1 = 426713070.440696 lpscbe1 = 1490.6611489301 wpscbe1 = 488.871169975975 ppscbe1 = -0.0019522282760703
+ pscbe2 = 4.17523356151092e-09 lpscbe2 = 2.14204712070922e-14 wpscbe2 = 1.02994388181522e-14 ppscbe2 = -4.13195473728039e-20
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 9.18114142186181e-11 lalpha0 = -1.13221159913114e-16 walpha0 = -1.20249283643804e-16 palpha0 = 1.48290531071154e-22
+ alpha1 = -3.85189284509951e-12 lalpha1 = 3.07916781804902e-17 walpha1 = 5.04498660910489e-18 palpha1 = -4.03291603218072e-23
+ beta0 = -29.498457816076 lbeta0 = -0.000232316440209147 wbeta0 = 7.79276410366345e-05 pbeta0 = 3.04274645495696e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -1.76249913515058e-10 lagidl = 9.54324750438669e-16 wagidl = 4.08908249577133e-16 pagidl = -1.13734698102165e-21
+ bgidl = 4070404912.6728 lbgidl = -12261.164613163 wbgidl = -4021.43888521489 pbgidl = 0.0160589647150062
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = 0.215767293164757 lkt1 = -2.55726900436609e-06 wkt1 = -1.10747457529843e-06 pkt1 = 4.2307613702025e-12
+ kt2 = 0.0276522015489231 lkt2 = -6.46848019459088e-07 wkt2 = -1.38616995657157e-07 pkt2 = 1.11625375620341e-12
+ at = 700484.210779479 lat = -2.73227595376442 wat = -0.963547626469386 pat = 4.05171332355793e-6
+ ute = 7.40343573436436 lute = -3.13336019634556e-05 wute = -1.29015561077682e-05 pute = 5.34713278751395e-11
+ ua1 = 1.70386756795036e-08 lua1 = -5.58201541001395e-14 wua1 = -2.54964267674012e-14 pua1 = 9.58494170733675e-20
+ ub1 = -9.13700837332206e-18 lub1 = 3.40385016447918e-23 wub1 = 1.45887910425019e-23 pub1 = -6.03621709381733e-29
+ uc1 = 1.20714519046778e-09 luc1 = -6.01616356044138e-15 wuc1 = -1.45499507151844e-15 puc1 = 6.95782790081299e-21
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.57 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 1.26e-06 wmax = 1.65e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.004443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.13309937680618+0*(0.005856/sqrt(l*w*mult))} lvth0 = 6.52865300238187e-08 wvth0 = 1.6281781663063e-07 pvth0 = -5.68750170316811e-14
+ k1 = 0.262056531028444 lk1 = 8.4849041147321e-07 wk1 = 2.30858618970434e-07 pk1 = -1.05147307192248e-12
+ k2 = 0.0957324515871884 lk2 = -3.29346412151091e-07 wk2 = -1.07936664382282e-07 pk2 = 4.15447174246221e-13
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 44830.6131584935 lvsat = -0.233251247530985 wvsat = -0.0166873716784494 pvsat = 3.61233080581679e-7
+ ua = 3.09892228816686e-09 lua = -6.28039116663418e-15 wua = -4.88441342057092e-15 pua = 7.19922120795389e-21
+ ub = -6.0803066611114e-19 lub = 2.01334461522432e-24 wub = 2.27472612323588e-24 pub = -1.85534352665691e-30
+ uc = -2.4633154526909e-10 luc = 2.32055286209232e-16 wuc = 2.38706309275638e-16 puc = -2.54211287877633e-22
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0281504448662749 lu0 = -3.37531846855121e-08 wu0 = -2.31358388506404e-08 pu0 = 4.06444856873366e-14
+ a0 = 1.4963528413622 la0 = -2.39939239784484e-06 wa0 = -3.68262177357714e-07 pa0 = 2.9312285082026e-12
+ keta = -0.0274058270029605 lketa = -1.02416663508307e-07 wketa = 5.06059054789188e-08 pketa = 9.22459795292096e-14
+ a1 = 0.0
+ a2 = 0.8
+ ags = -0.434971147811929 lags = 3.46225186172174e-06 wags = 8.73473338437298e-07 pags = -4.15799813437665e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.345784949781473+0*(0.0/sqrt(l*w*mult))} lvoff = 1.15822147745914e-08 wvoff = 8.59412474605751e-08 pvoff = -1.86455726124082e-14
+ nfactor = {0.211017464811619+0*(0.1/sqrt(l*w*mult))} lnfactor = 2.95024475308949e-06 wnfactor = 2.85505889272422e-06 pnfactor = -5.47670472384933e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = -0.18609657993379 leta0 = 1.06261358431964e-06 weta0 = 4.52295586189136e-07 peta0 = -1.80616915156135e-12
+ etab = 0.162625307030371 letab = -9.28951478326047e-07 wetab = -3.95403051147478e-07 petab = 1.57897802946317e-12
+ dsub = -0.444138037485999 ldsub = 4.00986258233826e-06 wdsub = 1.70677579694013e-06 pdsub = -6.81573264740132e-12
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.70974964528105 lpclm = -4.14761081481598e-06 wpclm = -3.90955810702429e-06 ppclm = 7.0706061973012e-12
+ pdiblc1 = 0.39
+ pdiblc2 = -0.00530281481429438 lpdiblc2 = 1.09988699462959e-08 wpdiblc2 = 9.37886269164132e-09 ppdiblc2 = -1.86952434000309e-14
+ pdiblcb = 0.543878313301866 lpdiblcb = 4.10452664097085e-07 wpdiblcb = -1.00703237359627e-06 ppdiblcb = -5.37587175270378e-13
+ drout = 0.56
+ pscbe1 = 800000134.108803 lpscbe1 = -0.000267324172455119 wpscbe1 = -0.000227950391490594 ppscbe1 = 4.54382177716983e-10
+ pscbe2 = 1.11778463431706e-08 lpscbe2 = -6.54332851319534e-15 wpscbe2 = -2.02310004718823e-15 ppscbe2 = 7.888515334637e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -8.21584610756616e-11 lalpha0 = 5.81499353954794e-16 walpha0 = 1.03626318588601e-16 palpha0 = -7.45720418596394e-22
+ alpha1 = -4.26684481638701e-10 lalpha1 = 1.71930512264835e-15 walpha1 = 5.58850488434739e-16 palpha1 = -2.25186171537118e-21
+ beta0 = -193.323014968594 lbeta0 = 0.000421890389201177 wbeta0 = 0.000327740822051358 pbeta0 = -6.93313823151279e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 2.66332297459237e-10 lagidl = -8.13055610769002e-16 wagidl = -2.61234337994005e-16 pagidl = 1.5387588793445e-21
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.362519145179734 lkt1 = -2.47975795240377e-07 wkt1 = -1.16702132407964e-07 pkt1 = 2.74272124655165e-13
+ kt2 = -0.176477384525888 lkt2 = 1.68310413537728e-07 wkt2 = 2.20638915650107e-07 pkt2 = -3.1837652614452e-13
+ at = -60799.1601499153 lat = 0.307785860136025 wat = 0.214427598618021 pat = -6.52339905842163e-7
+ ute = 0.667952381135571 lute = -4.43654034063966e-06 wute = 1.1047593901243e-07 pute = 1.50988584551249e-12
+ ua1 = 6.36131383769795e-09 lua1 = -1.31818393175071e-14 wua1 = -3.11156594048633e-15 pua1 = 6.45910170853693e-21
+ ub1 = -1.39515228047283e-18 lub1 = 3.12265351868547e-24 wub1 = -1.80307999769919e-24 pub1 = 5.09611057776103e-30
+ uc1 = -4.34624422706946e-10 luc1 = 5.39977423094566e-16 wuc1 = 2.79277610696139e-16 puc1 = 3.22908965635936e-23
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.58 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 1.26e-06 wmax = 1.65e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.004443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.17820063689786+0*(0.005856/sqrt(l*w*mult))} lvth0 = 1.55188585612456e-07 wvth0 = 2.24520873372474e-07 pvth0 = -1.79870064751356e-13
+ k1 = 0.802645567049158 lk1 = -2.29086256410248e-07 wk1 = -4.37237405411771e-07 pk1 = 2.80268121127493e-13
+ k2 = -0.11509478885164 lk2 = 9.09035376507616e-08 wk2 = 1.5661704056752e-07 pk2 = -1.11897778871007e-13
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -390963.785139197 lvsat = 0.635434286782936 wvsat = 0.614091071646121 pvsat = -8.96121560078033e-7
+ ua = 3.29318691110069e-09 lua = -6.66762622158385e-15 wua = -6.01703155420386e-15 pua = 9.45691197321352e-21
+ ub = -1.65175280460187e-18 lub = 4.09383561531915e-24 wub = 4.32573104914663e-24 pub = -5.94368958366198e-30
+ uc = -2.91060830445357e-10 luc = 3.21215870063922e-16 wuc = 3.26979210259922e-16 puc = -4.30169015779845e-22
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0236734912505302 lu0 = -2.48291029190109e-08 wu0 = -1.964468793724e-08 pu0 = 3.36854419079208e-14
+ a0 = -1.88878507956812 la0 = 4.34833165518654e-06 wa0 = 4.61032536682835e-06 pa0 = -6.99277922995015e-12
+ keta = -0.249028955554392 lketa = 3.39353140312146e-07 wketa = 3.62826382566213e-07 pketa = -5.30114961827023e-13
+ a1 = 0.0
+ a2 = 0.8
+ ags = 3.67528159780154 lags = -4.7308711257139e-06 wags = -5.32897519735221e-06 pags = 8.20557822505693e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.269419496643836+0*(0.0/sqrt(l*w*mult))} lvoff = -1.40639944851877e-07 wvoff = -2.52146264524148e-08 pvoff = 2.02925654781564e-13
+ nfactor = {3.38072621933057+0*(0.1/sqrt(l*w*mult))} lnfactor = -3.36805615622581e-06 wnfactor = -2.46675349428202e-06 pnfactor = 5.13146613604091e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = -1.16281092259415 leta0 = 3.00953539868956e-06 weta0 = 1.42020657959414e-06 peta0 = -3.7355429153333e-12
+ etab = 97.9650200521429 letab = -0.000195882181414759 wetab = -0.000128301119152594 petab = 2.56538302351689e-10
+ dsub = 3.867059549944 ldsub = -4.58381139419427e-06 wdsub = -5.11462311971374e-06 pdsub = 6.78162102632368e-12
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.221754719860793 lpclm = 1.69586823338714e-06 wpclm = 7.27012042452521e-07 ppclm = -2.1716452713166e-12
+ pdiblc1 = 0.42428281429169 lpdiblc1 = -6.83372364745678e-08 wpdiblc1 = -3.48048873590841e-08 ppdiblc1 = 6.93779045585817e-14
+ pdiblc2 = -0.000715794823729934 lpdiblc2 = 1.85538869234418e-09 wpdiblc2 = 1.21910126018066e-09 ppdiblc2 = -2.43008086776599e-15
+ pdiblcb = 1.41455173436522 lpdiblcb = -1.3250937516985e-06 wpdiblcb = -2.40759343507404e-06 ppdiblcb = 2.25420440989358e-12
+ drout = 0.868453341004798 ldrout = -6.14851765851821e-07 wdrout = -8.60980115275817e-07 pdrout = 1.71622438102367e-12
+ pscbe1 = 800000000.0
+ pscbe2 = 1.18969441836019e-08 lpscbe2 = -7.97673356424496e-15 wpscbe2 = -2.05491499482408e-15 ppscbe2 = 7.95193327872753e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.18395971471157e-10 lalpha0 = -2.16941017509216e-16 walpha0 = -5.3915813995363e-16 palpha0 = 5.35566268425259e-22
+ alpha1 = 7.69444931387629e-10 lalpha1 = -6.64985089254725e-16 walpha1 = -1.13788380045566e-15 palpha1 = 1.13030321857702e-21
+ beta0 = 27.7942051024633 lbeta0 = -1.88709680208248e-05 wbeta0 = -4.01513503565217e-05 pbeta0 = 4.00196240118995e-11
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -3.81499121616201e-10 lagidl = 4.78291374467994e-16 wagidl = 1.01803054651621e-15 pagidl = -1.01124842701532e-21
+ bgidl = 140972920.602244 lbgidl = 1712.33132039256 wbgidl = 1125.10401682999 pbgidl = -0.00224271259069986
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.738360763569044 lkt1 = 5.01203584676532e-07 wkt1 = 4.05996308599238e-07 pkt1 = -7.67642540345248e-13
+ kt2 = -0.179245092622563 lkt2 = 1.73827391259737e-07 wkt2 = 1.99002595075393e-07 pkt2 = -2.75248026162759e-13
+ at = -17354.309577376 lat = 0.221185588585461 wat = 0.0123462150321751 pat = -2.4952340484792e-7
+ ute = -5.3249347975136 lute = 7.50930940227453e-06 wute = 6.19020637415626e-06 pute = -1.06090718606162e-11
+ ua1 = -2.39547311000422e-09 lua1 = 4.2733968632517e-15 wua1 = 3.0500424111103e-15 pua1 = -5.82306635981799e-21
+ ub1 = -2.76214515581494e-19 lub1 = 8.92232352292501e-25 wub1 = 1.68681372123368e-24 pub1 = -1.86042718814917e-30
+ uc1 = -5.77073994705279e-10 luc1 = 8.2392756804258e-16 wuc1 = 8.55619595892063e-16 puc1 = -1.11655348352288e-21
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.59 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 1.26e-06 wmax = 1.65e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.004443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.01004200544915+0*(0.005856/sqrt(l*w*mult))} lvth0 = -1.18497730335388e-08 wvth0 = -1.55089902675302e-08 pvth0 = 5.85607199370768e-14
+ k1 = 0.885348114424805 lk1 = -3.11237839415278e-07 wk1 = -6.37192030645503e-07 pk1 = 4.78890648647919e-13
+ k2 = -0.146932329533757 lk2 = 1.22528976636855e-07 wk2 = 2.24390840157271e-07 pk2 = -1.79220069407891e-13
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 346418.317349862 lvsat = -0.0970353761393405 wvsat = -0.470515839931597 pvsat = 1.81259700254754e-7
+ ua = -5.38320252327834e-09 lua = 1.95096110638335e-15 wua = 6.5723794001045e-15 pua = -3.04862832531725e-21
+ ub = 3.54116292643623e-18 lub = -1.06448491111878e-24 wub = -3.34145336545218e-24 pub = 1.67241604836677e-30
+ uc = 2.27378112630769e-11 luc = 9.50775490654963e-18 wuc = -1.28278950348005e-16 puc = 2.2056214962113e-23
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = -0.0105184400572399 lu0 = 9.13504174238687e-09 wu0 = 2.91537287745804e-08 pu0 = -1.47878797517655e-14
+ a0 = 4.3839777211127 la0 = -1.88264199971615e-06 wa0 = -5.55964943632238e-06 pa0 = 3.10944320106198e-12
+ keta = 0.126745361892265 lketa = -3.39177686316813e-08 wketa = -2.21360021383582e-07 pketa = 5.0179592299658e-14
+ a1 = 0.0
+ a2 = 0.622863910459608 la2 = 1.75956008911874e-07 wa2 = 2.32002611614032e-07 pa2 = -2.30457010215458e-13
+ ags = -2.12186353869076 lags = 1.02765342987908e-06 wags = 4.07772071829569e-06 pags = -1.13845028240093e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.359410493563707+0*(0.0/sqrt(l*w*mult))} lvoff = -5.12484679534861e-08 wvoff = 1.47025668625934e-07 pvoff = 3.18328245490271e-14
+ nfactor = {-0.988608471007618+0*(0.1/sqrt(l*w*mult))} lnfactor = 9.72170026405347e-07 wnfactor = 3.81650243684772e-06 pnfactor = -1.10993074407564e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 3.22547100492347 leta0 = -1.34951179462693e-06 weta0 = -4.64959550394482e-06 peta0 = 2.29382214672513e-12
+ etab = -197.137625864247 letab = 9.72544906745357e-05 wetab = 0.000258181261645271 petab = -1.27369332825301e-10
+ dsub = -1.67741657416397 ldsub = 9.23727429974888e-07 wdsub = 3.24392486851004e-06 pdsub = -1.52124231520255e-12
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.347851242867 lpclm = -8.5661901441696e-07 wpclm = -2.91801340946853e-06 ppclm = 1.44909702104375e-12
+ pdiblc1 = 0.407050002259573 lpdiblc1 = -5.12192294362095e-08 wpdiblc1 = 2.60967824871713e-07 ppdiblc1 = -2.24424369863334e-13
+ pdiblc2 = 0.00152615705793975 lpdiblc2 = -3.71627305889825e-10 wpdiblc2 = -2.12718248138569e-09 ppdiblc2 = 8.93909931514041e-16
+ pdiblcb = 1.04478401132076 lpdiblcb = -9.57789421224963e-07 wpdiblcb = -1.40114126451208e-06 ppdiblcb = 1.25445722369191e-12
+ drout = -0.491044122009595 ldrout = 7.3558872506397e-07 wdrout = 1.72196023055163e-06 pdrout = -8.49508416219882e-13
+ pscbe1 = 800000000.0
+ pscbe2 = -1.5373240883963e-09 lpscbe2 = 5.36803561252522e-15 wpscbe2 = 1.1855759218561e-14 ppscbe2 = -5.86606802304801e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 7.04102368697252 lbeta0 = 1.743955700076e-06 wbeta0 = 2.26701701300324e-06 pbeta0 = -2.11615219420968e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 5.59851478234573e-10 lagidl = -4.56787947686574e-16 wagidl = -9.62015589866671e-16 pagidl = 9.5560664200698e-22
+ bgidl = 2718054158.79551 lbgidl = -847.58140259186 wbgidl = -2250.20803365998 pbgidl = 0.00111011313090975
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = 0.0372088399887707 lkt1 = -2.69199174182381e-07 wkt1 = -7.28701958307797e-07 pkt1 = 3.59496366707652e-13
+ kt2 = 0.0460055339764513 lkt2 = -4.99226156648746e-08 wkt2 = -1.55142372751517e-07 pkt2 = 7.65376278884877e-14
+ at = 305573.687518636 lat = -0.0995910621938978 wat = -0.424504856285423 pat = 1.8441736463256e-7
+ ute = 5.00824121046288 lute = -2.75502698713682e-06 wute = -9.35388944844504e-06 pute = 4.8314691956149e-12
+ ua1 = 3.23896573225266e-09 lua1 = -1.32350534743806e-15 wua1 = -5.58668666250101e-15 pua1 = 2.75612482470492e-21
+ ub1 = 1.26843189565092e-18 lub1 = -6.42123624548278e-25 wub1 = -1.12526300402819e-24 pub1 = 9.32915481968996e-31
+ uc1 = 4.77400120260054e-10 luc1 = -2.23521640368855e-16 wuc1 = -5.33268050757295e-16 puc1 = 2.63081393624503e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.60 pmos
* DC IV MOS Parameters
+ lmin = 2.5e-07 lmax = 5e-07 wmin = 1.26e-06 wmax = 1.65e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.006443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.960607295430903+0*(0.007356/sqrt(l*w*mult))} lvth0 = -3.62377940045217e-08 wvth0 = 1.53457138600076e-08 pvth0 = 4.33389219122074e-14
+ k1 = -0.870839999532857 lk1 = 5.55156492348367e-07 wk1 = 1.71670363862158e-06 pk1 = -6.82375533036964e-13
+ k2 = 0.496158449118115 lk2 = -1.94732141921703e-07 wk2 = -6.43213045632426e-07 pk2 = 2.48801896399827e-13
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 202824.348665743 lvsat = -0.0261950148166546 wvsat = -0.225333536452963 pvsat = 6.03019530212122e-8
+ ua = 2.99483138063512e-10 lua = -8.52523672411721e-16 wua = -1.33540609511111e-15 pua = 8.52582755321427e-22
+ ub = 6.31707987743998e-19 lub = 3.7085976942577e-25 wub = 6.97421314009498e-25 pub = -3.20114308249495e-31
+ uc = 1.1037409937167e-10 luc = -3.37265561963678e-17 wuc = -2.00968368565343e-16 puc = 5.79166671666178e-23
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.015263691195774 lu0 = -3.58426332571251e-09 wu0 = -8.00502537772731e-09 pu0 = 3.54394570422566e-15
+ a0 = 1.65025854981243 la0 = -5.33994451185211e-07 wa0 = -2.62447342981096e-07 pa0 = 4.96132114737178e-13
+ keta = 0.408858957758571 lketa = -1.73095125789173e-07 wketa = -6.0900329893816e-07 pketa = 2.41418751561879e-13
+ a1 = 0.0
+ a2 = 0.251172969660389 la2 = 3.5932527426388e-07 wa2 = 1.07103061381042e-06 pa2 = -6.44381406763023e-13
+ ags = -2.53523781434261 lags = 1.23158666828061e-06 wags = 6.17546614783037e-06 pags = -2.17334781711671e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.521949906309723+0*(0.0/sqrt(l*w*mult))} lvoff = 2.89384008518076e-08 wvoff = 4.41891599783223e-07 pvoff = -1.13635744196248e-13
+ nfactor = {0.282152463094171+0*(0.1/sqrt(l*w*mult))} lnfactor = 3.45255368697438e-07 wnfactor = 1.40698415489704e-06 pnfactor = 7.877618610534e-14
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 1.32617658651253 leta0 = -4.1251768483692e-07 weta0 = -1.09517576200741e-06 peta0 = 5.40291820077214e-13
+ etab = -0.00395776844010065 letab = 9.61123486551509e-10 wetab = 5.2471802157573e-09 petab = -1.29420113966165e-15
+ dsub = 0.308547421412642 ldsub = -5.60240756748854e-08 wdsub = -3.84323373835187e-07 pdsub = 2.68710416179558e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.31250524601823 lpclm = 4.558359350967e-07 wpclm = 1.21556787285796e-06 ppclm = -5.90155701616637e-13
+ pdiblc1 = 0.465892152337624 lpdiblc1 = -8.02482980714149e-08 wpdiblc1 = -7.9810921112226e-07 ppdiblc1 = 2.98058576919861e-13
+ pdiblc2 = 0.00474571276608955 lpdiblc2 = -1.95995647983704e-09 wpdiblc2 = -1.89493752232203e-08 ppdiblc2 = 9.19293685438523e-15
+ pdiblcb = -1.97568158996172 lpdiblcb = 5.32321037580538e-07 wpdiblcb = 2.80985803510685e-06 ppdiblcb = -8.22988748783494e-13
+ drout = 0.898895496875351 ldrout = 4.98786933625088e-08 wdrout = 8.56938533734916e-07 pdrout = -4.22760342355716e-13
+ pscbe1 = 799767456.074087 lpscbe1 = 0.114722755322418 wpscbe1 = 0.395264724227673 ppscbe1 = -1.94999108521412e-7
+ pscbe2 = 9.40276673535493e-09 lpscbe2 = -2.91269142825731e-17 wpscbe2 = 2.48841346709769e-17 ppscbe2 = -2.94477709118472e-23
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 13.396648879577 lbeta0 = -1.39151572119309e-06 wbeta0 = -6.04980482296609e-06 pbeta0 = 1.98685205670376e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -1.12677109608235e-08 lagidl = 5.37819805087344e-15 wagidl = 1.5608228168974e-14 pagidl = -7.21912427349195e-21
+ bgidl = 1906629732.22925 lbgidl = -447.274898838516 wbgidl = -1541.03681564476 pbgidl = 0.000760252020556555
+ cgidl = 1314.81899247236 lcgidl = -0.000500648772108331 wcgidl = -0.00132915125980254 pcgidl = 6.55720824208464e-10
+ egidl = -5.2700921379826 legidl = 2.64927051516806e-06 wegidl = 7.03343629100403e-06 pegidl = -3.46986139293135e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.411109332528258 lkt1 = -4.80267835891742e-08 wkt1 = -1.22902104300533e-07 pkt1 = 6.06322783314164e-14
+ kt2 = 0.0917427465178488 lkt2 = -7.24865206256225e-08 wkt2 = -2.40370290969696e-07 pkt2 = 1.18583798606408e-13
+ at = 183751.546951822 lat = -0.0394915710109467 wat = -0.157517563693496 pat = 5.27023876798438e-8
+ ute = -0.470047706110753 lute = -5.23788896122136e-08 wute = 2.29902898210111e-07 pute = 1.03420246900739e-13
+ ua1 = 1.5568073272951e-09 lua1 = -4.93632684253113e-16 wua1 = -1.11461985279068e-15 pua1 = 5.49884328936051e-22
+ ub1 = -2.96320798163869e-19 lub1 = 1.29828339912921e-25 wub1 = 1.25387204457542e-24 pub1 = -2.40802244639012e-31
+ uc1 = 4.73155848733005e-11 luc1 = -1.13445958502243e-17 wuc1 = 1.5618346075442e-19 puc1 = -7.70512361616663e-26
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.24e-6
+ sbref = 1.24e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.61 pmos
* DC IV MOS Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 1.26e-06 wmax = 1.65e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.006443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.878886907244986+0*(0.007356/sqrt(l*w*mult))} lvth0 = -5.61234698249064e-08 wvth0 = 1.58236831312625e-07 pvth0 = 8.5680831735206e-15
+ k1 = 3.09060327611239 lk1 = -4.08813191460595e-07 wk1 = -5.06654607030933e-06 pk1 = 9.68246884634865e-13
+ k2 = -0.941669914875341 lk2 = 1.55146136515737e-07 wk2 = 1.83911630929196e-06 pk2 = -3.55243164168764e-13
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 70301.0671297982 lvsat = 0.00605293546573915 wvsat = 0.219363306565091 pvsat = -4.79096873651152e-8
+ ua = -5.60992647605409e-09 lua = 5.85460244268429e-16 wua = 7.49106940890682e-15 pua = -1.29523414087529e-21
+ ub = 3.80296353054249e-18 lub = -4.00827211847729e-25 wub = -4.49599295230153e-24 pub = 9.436407324861e-31
+ uc = -9.89370266206271e-11 luc = 1.7206794580346e-17 wuc = 1.29091223672635e-16 puc = -2.23993738893872e-23
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = -0.00607121728030889 lu0 = 1.60733063304055e-09 wu0 = 2.18615547004308e-08 pu0 = -3.72372815883316e-15
+ a0 = -2.46687383977989 la0 = 4.67860310233404e-07 wa0 = 3.4030841850462e-06 pa0 = -3.95830996229929e-13
+ keta = -1.08381757113888 lketa = 1.90129795399675e-07 wketa = 1.28616347147215e-06 pketa = -2.19747340016225e-13
+ a1 = 0.0
+ a2 = 4.4666105048153 la2 = -6.66450864665647e-07 wa2 = -5.69302234185812e-06 pa2 = 1.00156971136345e-12
+ ags = 5.68563527163015 lags = -7.68864146713827e-07 wags = -9.58031765194225e-06 pags = 1.66063310115236e-12
+ b0 = 0.0
+ b1 = 1.75247592434801e-23 lb1 = -4.26443986478995e-30 wb1 = -2.97875728309831e-29 pb1 = 7.24844839754578e-36
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.212808651804103+0*(0.0/sqrt(l*w*mult))} lvoff = -4.62874137370809e-08 wvoff = -9.6525924582703e-09 pvoff = -3.75788354458727e-15
+ nfactor = {3.03855510498472+0*(0.1/sqrt(l*w*mult))} lnfactor = -3.25482137374923e-07 wnfactor = -2.83630738169255e-06 pnfactor = 1.11133026203598e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = -1.48955334860311 leta0 = 2.72656406114251e-07 weta0 = 3.49637538648327e-06 peta0 = -5.77007053294212e-13
+ etab = 0.583180912759274 letab = -1.41912028919142e-07 wetab = -6.61760958351805e-07 petab = 1.61014225283092e-13
+ dsub = -0.419015932804587 ldsub = 1.21019735813627e-07 wdsub = 2.53407159296825e-06 pdsub = -4.41445978252457e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 3.78991247095034 lpclm = -5.42438187314997e-07 wpclm = -4.08034707481284e-06 ppclm = 6.98541649919682e-13
+ pdiblc1 = -0.212048977222925 lpdiblc1 = 8.47205405135901e-08 wpdiblc1 = 1.88722795190995e-06 ppdiblc1 = -3.55385997658071e-13
+ pdiblc2 = -0.0357092232155182 lpdiblc2 = 7.88426673205544e-09 wpdiblc2 = 8.96521533276172e-08 ppdiblc2 = -1.72339419001185e-14
+ pdiblcb = 0.114993147851663 lpdiblcb = 2.35804282305033e-08 wpdiblcb = -9.31792145159875e-07 ppdiblcb = 8.74969227822502e-14
+ drout = 1.36108751115946 ldrout = -6.25901870093584e-08 wdrout = -3.06049476333898e-06 pdrout = 5.30500041287652e-13
+ pscbe1 = 800830514.021122 lpscbe1 = -0.143959639392961 wpscbe1 = -1.4116597293887 ppscbe1 = 2.44694274172813e-7
+ pscbe2 = 8.06601424215027e-09 lpscbe2 = 2.96155763908869e-16 wpscbe2 = 9.18436028947751e-16 ppscbe2 = -2.46882901761371e-22
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 7.20416726554275 lbeta0 = 1.15350369802766e-07 wbeta0 = 4.36024234050139e-06 pbeta0 = -5.46307999960091e-13
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 3.52389060251324e-08 lagidl = -5.93862911325509e-15 wagidl = -4.60229080829501e-14 pagidl = 7.77807315977877e-21
+ bgidl = -2213402715.05922 lbgidl = 555.285556819766 wbgidl = 5461.95620038073 pbgidl = -0.000943842293977056
+ cgidl = -3324.35354454415 lcgidl = 0.000628238194704193 wcgidl = 0.00474696878500905 pcgidl = -8.22830075255898e-10
+ egidl = 19.278900492795 legidl = -3.32443225362009e-06 wegidl = -2.51194153250144e-05 pegidl = 4.35414921360734e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.967724069659923 lkt1 = 8.74187333149706e-08 wkt1 = 1.0054723644546e-06 pkt1 = -2.1394410814652e-13
+ kt2 = -0.398296571328263 lkt2 = 4.67586669004146e-08 wkt2 = 8.30760457021826e-07 pkt2 = -1.42063015348353e-13
+ at = -170851.234395878 lat = 0.0467967605966398 wat = 0.334981305312889 pat = -6.71413021064321e-8
+ ute = -0.942181992289765 lute = 6.2509323318015e-08 wute = 1.09154383237499e-06 pute = -1.06249734737074e-13
+ ua1 = -1.84132780195131e-09 lua1 = 3.33262721827451e-16 wua1 = 3.75631921824495e-15 pua1 = -6.35400242731618e-22
+ ub1 = 2.37210092666667e-19 wub1 = 2.64292757168557e-25
+ uc1 = 3.76355683135322e-12 luc1 = -7.46732450552953e-19 wuc1 = -5.37646616435935e-18 puc1 = 1.26925265831427e-24
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.62 pmos
* DC IV MOS Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 1.26e-06 wmax = 1.65e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.006443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.41151918892007+0*(0.007356/sqrt(l*w*mult))} lvth0 = 3.62019446160894e-08 wvth0 = 9.57093991088551e-07 pvth0 = -1.29904219187719e-13
+ k1 = -2.26758269068731 lk1 = 5.19964047652529e-07 wk1 = 3.28050999080543e-06 pk1 = -4.78615118886645e-13
+ k2 = 1.270846046865 lk2 = -2.2836695526041e-07 wk2 = -1.52134750859296e-06 pk2 = 2.27252913095773e-13
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 609409.86501181 lvsat = -0.0873951053415329 wvsat = -0.679172091022197 pvsat = 1.0784064138187e-7
+ ua = 1.51832618172493e-10 lua = -4.13271553606618e-16 wua = -1.68589330927599e-15 pua = 2.95482222769081e-22
+ ub = -1.92628253230173e-18 lub = 5.9226884219356e-25 wub = 3.72979820356283e-24 pub = -4.82201454889115e-31
+ uc = 2.58967002538763e-12 luc = -3.91639962880931e-19 wuc = -2.66739034501011e-18 puc = 4.39400747203288e-25
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0106864132997624 lu0 = -1.29740353644785e-09 wu0 = -7.35355871177798e-09 pu0 = 1.34036116981227e-15
+ a0 = -0.855173815380581 la0 = 1.88491451404077e-07 wa0 = 3.63354841529781e-06 pa0 = -4.35779204973282e-13
+ keta = -0.832689077893654 lketa = 1.46599684637534e-07 wketa = 1.42392918628321e-06 pketa = -2.43627373490145e-13
+ a1 = 0.0
+ a2 = -3.2019090525702 la2 = 6.62794978372442e-07 wa2 = 3.92372605858992e-06 pa2 = -6.6537822287341e-13
+ ags = 1.25
+ b0 = 0.0
+ b1 = -4.08911049014536e-23 lb1 = 5.86124919436455e-30 wb1 = 6.95043366056275e-29 pb1 = -9.96261260037743e-36
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.325624990069805+0*(0.0/sqrt(l*w*mult))} lvoff = -2.67320552947812e-08 wvoff = -3.46911122829019e-07 pvoff = 5.47018355928172e-14
+ nfactor = {-18.7383369998885+0*(0.1/sqrt(l*w*mult))} lnfactor = 3.44928078629959e-06 wnfactor = 2.51646927990893e-05 pnfactor = -3.74230710730038e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = -2.40631671785476 leta0 = 4.31566335013593e-07 weta0 = 3.43301549625914e-06 peta0 = -5.66024376642542e-13
+ etab = -0.861273939966609 letab = 1.08466886342657e-07 wetab = 9.81422155772066e-07 petab = -1.23811849352912e-13
+ dsub = 0.37068240177151 ldsub = -1.58649941051246e-08 wdsub = -7.31692156842309e-08 pdsub = 1.04879290377462e-14
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 3.71046415834999 lpclm = -5.28666775705477e-07 wpclm = -4.00898575898727e-06 ppclm = 6.86172022157109e-13
+ pdiblc1 = 3.47367782170907 lpdiblc1 = -5.54155971359683e-07 wpdiblc1 = -4.28707368099367e-06 ppdiblc1 = 7.14855098786177e-13
+ pdiblc2 = 0.0900650406287515 lpdiblc2 = -1.39171926141826e-08 wpdiblc2 = -1.17032870312573e-07 ppdiblc2 = 1.85924267276248e-14
+ pdiblcb = -0.986217486520106 lpdiblcb = 2.14462077171237e-07 wpdiblcb = 1.6746124030252e-06 ppdiblcb = -3.64292028791054e-13
+ drout = 1.0
+ pscbe1 = 800000000.0
+ pscbe2 = 9.62513689678327e-09 lpscbe2 = 2.59005612000915e-17 wpscbe2 = 1.00109926457981e-15 ppscbe2 = -2.6121158169936e-22
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 15.8812623700667 lbeta0 = -1.3887199414252e-06 wbeta0 = -3.93890592882478e-06 pbeta0 = 8.92249762748357e-13
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 6.21001594322295e-09 lagidl = -9.06819364237071e-16 wagidl = -9.88484558059839e-15 pagidl = 1.51397368174612e-21
+ bgidl = 942691899.894409 lbgidl = 8.21442845293495 wbgidl = 97.4089961512946 pbgidl = -1.39624106903343e-5
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = 0.713698580275306 lkt1 = -2.04035705979502e-07 wkt1 = -1.32191798122296e-06 pkt1 = 1.89481079592537e-13
+ kt2 = -0.169356806016125 lkt2 = 7.07470586073925e-09 wkt2 = 6.46446916965319e-08 pkt2 = -9.26604081839745e-15
+ at = 573319.148647231 lat = -0.0821962452592865 wat = -0.622109915146003 pat = 9.87589758654713e-8
+ ute = -2.34524425071694 lute = 3.05713329069265e-07 wute = 2.76520966930472e-06 pute = -3.96359623578799e-13
+ ua1 = -2.37427591297519e-11 lua1 = 1.82061656748483e-17 wua1 = 2.46448790969746e-17 pua1 = 1.14407238676131e-23
+ ub1 = -3.92043284578177e-19 lub1 = 1.09073521904867e-25 wub1 = 1.52706593140277e-24 pub1 = -2.18886576475411e-31
+ uc1 = -3.3955526523995e-11 luc1 = 5.79141802009639e-18 wuc1 = 1.12435588772182e-17 puc1 = -1.61162924234271e-24
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.63 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 1e-06 wmax = 1.26e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.004443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.0053647+0*(0.005856/sqrt(l*w*mult))}
+ k1 = 0.49177002
+ k2 = -0.002473247
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 55237.817
+ ua = -1.3943119e-9
+ ub = 1.565972e-18
+ uc = -3.8916596e-11
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0072382252
+ a0 = 1.248405
+ keta = 0.0066402373
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.25185017
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.29956891+0*(0.0/sqrt(l*w*mult))}
+ nfactor = {1.7720538+0*(0.1/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.0017402344
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00056783834
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 799985290.0
+ pscbe2 = 1.0771971e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.0
+ alpha1 = 0.0
+ beta0 = 30.0
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.4670794e-10
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.54561
+ kt2 = -0.052484
+ at = 10000.0
+ ute = -1.2595
+ ua1 = -2.5605e-10
+ ub1 = 4.9434e-19
+ uc1 = 8.1951e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.64 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 1e-06 wmax = 1.26e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.004443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.0053647+0*(0.005856/sqrt(l*w*mult))}
+ k1 = 0.49177002
+ k2 = -0.002473247
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 55237.817
+ ua = -1.3943119e-9
+ ub = 1.565972e-18
+ uc = -3.8916596e-11
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0072382252
+ a0 = 1.248405
+ keta = 0.0066402373
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.25185017
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.29956891+0*(0.0/sqrt(l*w*mult))}
+ nfactor = {1.7720538+0*(0.1/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.0017402344
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00056783834
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 799985290.0
+ pscbe2 = 1.0771971e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.0
+ alpha1 = 0.0
+ beta0 = 30.0
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.4670794e-10
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.54561
+ kt2 = -0.052484
+ at = 10000.0
+ ute = -1.2595
+ ua1 = -2.5605e-10
+ ub1 = 4.9434e-19
+ uc1 = 8.1951e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.65 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 1e-06 wmax = 1.26e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.004443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.0074140810616+0*(0.005856/sqrt(l*w*mult))} lvth0 = 1.63813955161699e-8
+ k1 = 0.533711539863405 lk1 = -3.35252744501912e-7
+ k2 = -0.015204835164966 lk2 = 1.01767887479373e-07 wk2 = 3.30872245021211e-24
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 67709.0584957215 lvsat = -0.0996868485549278
+ ua = -1.96104979334727e-09 lua = 4.53012753893265e-15
+ ub = 1.85327925148432e-18 lub = -2.29654397096517e-24
+ uc = -2.32886427786375e-11 luc = -1.24919512346539e-16
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0046760248637794 lu0 = 2.0480533311125e-8
+ a0 = 1.3219165622399 la0 = -5.87602763891554e-7
+ keta = 0.0100523898791525 lketa = -2.72744888727377e-8
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.199837851034395 lags = 4.15752045655893e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.318274014675695+0*(0.0/sqrt(l*w*mult))} lvoff = 1.49516223998211e-7
+ nfactor = {1.4620747314211+0*(0.1/sqrt(l*w*mult))} lnfactor = 2.47776746807634e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.0344627685079662 lpclm = 2.89382838858357e-07 wpclm = -9.92616735063633e-24 ppclm = -2.52435489670724e-29
+ pdiblc1 = 0.39
+ pdiblc2 = 9.85732448773808e-05 lpdiblc2 = 3.75099451691726e-9
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 799970624.466194 lpscbe1 = 0.117226568654587
+ pscbe2 = 1.20389481292726e-08 lpscbe2 = -1.01273764325456e-14
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.0
+ alpha1 = 0.0
+ beta0 = 30.0
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.35955228517575e-10 lagidl = 8.59500572955045e-17
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.629799548385 lkt1 = 6.72955516308661e-7
+ kt2 = -0.0781831266990001 lkt2 = 2.05421806009931e-7
+ at = -35193.10531325 lat = 0.361243766038403 wat = 1.38777878078145e-17 pat = -5.29395592033938e-23
+ ute = -2.44701888775 lute = 9.49223985116981e-6
+ ua1 = -2.428076454925e-09 lua1 = 1.73617415991573e-14 wua1 = 7.88860905221012e-31
+ ub1 = 2.00166536148e-18 lub1 = -1.20485610902818e-23
+ uc1 = 9.624331106095e-11 luc1 = -7.03799111305513e-16 wuc1 = -2.46519032881566e-32 puc1 = -2.82118644197349e-37
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.66 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 1e-06 wmax = 1.26e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.004443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.0087865031501+0*(0.005856/sqrt(l*w*mult))} lvth0 = 2.18619407942096e-8
+ k1 = 0.438319171852289 lk1 = 4.56812235868604e-8
+ k2 = 0.01332183338898 lk2 = -1.21487420705046e-8
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 32089.65415263 lvsat = 0.0425534723457048
+ ua = -6.30371477103069e-10 lua = -7.83720747101319e-16
+ ub = 1.12874327553622e-18 lub = 5.96773074155461e-25
+ uc = -6.4077122012637e-11 luc = 3.79626717408017e-17
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0104860229284 lu0 = -2.72075274025099e-9
+ a0 = 1.2151813426064 la0 = -1.61372955390757e-7
+ keta = 0.0112322389301054 lketa = -3.19860249221719e-08 pketa = 1.26217744835362e-29
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.231933635768609 lags = 2.87582728836931e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.28016803107749+0*(0.0/sqrt(l*w*mult))} lvoff = -2.65384833187796e-9
+ nfactor = {2.3908807178428+0*(0.1/sqrt(l*w*mult))} lnfactor = -1.23126877212893e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.1592351855 leta0 = -3.16412877194199e-7
+ etab = -0.139268494014963 letab = 2.76612509352725e-7
+ dsub = 0.8590007 ldsub = -1.1940108573366e-6
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.275233282675524 lpclm = 1.2508608823632e-06 ppclm = -2.01948391736579e-28
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0018580315657347 lpdiblc2 = -3.27511725517847e-9
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 799999960.066619 lpscbe1 = 7.96007225289941e-5
+ pscbe2 = 9.63319118340849e-09 lpscbe2 = -5.20375801862541e-16
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -3.038830824303e-12 lalpha0 = 1.21350786062605e-17
+ alpha1 = 2.9141211206745e-15 lalpha1 = -1.16370706077921e-20
+ beta0 = 56.9100629999999 lbeta0 = -0.000107460977160294
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 6.68775207909697e-11 lagidl = 3.6180069251305e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.451622277389999 lkt1 = -3.85665506919725e-8
+ kt2 = -0.00801757949699999 lkt2 = -7.4772939922609e-8
+ at = 102918.248221 lat = -0.190281550261352
+ ute = 0.75230175845 lute = -3.28372885948521e-06 wute = 4.2351647362715e-22 pute = -1.41363874215605e-27
+ ua1 = 3.98560513679e-09 lua1 = -8.25025682093871e-15
+ ub1 = -2.77182014511e-18 lub1 = 7.01357997563328e-24 pub1 = -2.80259692864963e-45
+ uc1 = -2.21393444354e-10 luc1 = 5.64631814289714e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.67 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 1e-06 wmax = 1.26e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.004443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.006776922084+0*(0.005856/sqrt(l*w*mult))} lvth0 = 1.78561664910749e-8
+ k1 = 0.468810858652519 lk1 = -1.50990143961379e-8
+ k2 = 0.00448373627148799 lk2 = 5.46857276148265e-9
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 77900.294865342 lvsat = -0.0487626185912911
+ ua = -1.30087102961762e-09 lua = 5.52811489908928e-16
+ ub = 1.65098192376424e-18 lub = -4.44225068426082e-25
+ uc = -4.14092499588139e-11 luc = -7.22205900322166e-18
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.00867459456899998 lu0 = 8.90036242818672e-10
+ a0 = 1.6312399809578 la0 = -9.90718449444858e-7
+ keta = 0.0279922647790546 lketa = -6.53944213278645e-08 wketa = 6.61744490042422e-24 pketa = 2.52435489670724e-29
+ a1 = 0.0
+ a2 = 0.8
+ ags = -0.393439099563341 lags = 1.53416196633805e-6
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.2886710916924+0*(0.0/sqrt(l*w*mult))} lvoff = 1.42956255081255e-8
+ nfactor = {1.4973376453944+0*(0.1/sqrt(l*w*mult))} lnfactor = 5.4986458881922e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = -0.078470371 leta0 = 1.57414641388398e-07 weta0 = 2.31610571514848e-23 peta0 = 3.39210189245035e-29
+ etab = 0.00595669402992639 letab = -1.2870376534299e-08 petab = 4.73316543132607e-30
+ dsub = -0.0380014000000002 ldsub = 5.940175146732e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.333325541317719 lpclm = 3.77974532621591e-8
+ pdiblc1 = 0.39770896841646 lpdiblc1 = -1.536657968533e-8
+ pdiblc2 = 0.000215
+ pdiblcb = -0.4236676 lpdiblcb = 3.960116764488e-7
+ drout = 0.2110872461536 ldrout = 6.95501050926675e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 1.032799802395e-08 lpscbe2 = -1.90536067977383e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -9.32561383513941e-11 lalpha0 = 1.91968665957697e-16 walpha0 = 6.16297582203915e-33 palpha0 = -4.11423022787801e-38
+ alpha1 = -9.93396282422415e-11 lalpha1 = 1.98011627638892e-16 walpha1 = -4.42301848790681e-32 palpha1 = 5.21396029436995e-38
+ beta0 = -2.86171356345561 lbeta0 = 1.16843763911515e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 3.9577639605148e-10 lagidl = -2.93805933700985e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.428378914775259 lkt1 = -8.48984286397128e-8
+ kt2 = -0.0273048137834199 lkt2 = -3.63269629045852e-8
+ at = -7927.86288261802 lat = 0.030672215153712 pat = -1.32348898008484e-23
+ ute = -0.598656317553001 lute = -5.90812790181536e-7
+ ua1 = -6.673817948866e-11 lua1 = -1.72566899554433e-16
+ ub1 = 1.01168299679436e-18 lub1 = -5.28220610244075e-25
+ uc1 = 7.6199295177312e-11 luc1 = -2.85711019421528e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.68 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 1e-06 wmax = 1.26e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.004443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.021883259604+0*(0.005856/sqrt(l*w*mult))} lvth0 = 3.28618655905177e-8
+ k1 = 0.398846243563881 lk1 = 5.43994964267828e-8
+ k2 = 0.0243921037457624 lk2 = -1.43071651686781e-08 wk2 = 1.32348898008484e-23
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -12824.776391484 lvsat = 0.041358042240822
+ ua = -3.6513148601276e-10 lua = -3.76694156856437e-16
+ ub = 9.89933100099282e-19 lub = 2.12419847975621e-25
+ uc = -7.52043260124921e-11 luc = 2.63478742537868e-17
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0117406951944 lu0 = -2.1556380202149e-9
+ a0 = 0.139135158719601 la0 = 4.9144597046759e-7
+ keta = -0.0422650138775481 lketa = 4.39480333832778e-9
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.991513061907201 lags = 1.58436356167227e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.24715506755244+0*(0.0/sqrt(l*w*mult))} lvoff = -2.69438188790144e-8
+ nfactor = {1.92532561224+0*(0.1/sqrt(l*w*mult))} lnfactor = 1.24727877808744e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = -0.32453716 leta0 = 4.0184213344008e-7
+ etab = -0.013900565275 letab = 6.85459370913795e-9
+ dsub = 0.799349363827521 ldsub = -2.37754818365702e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.11992164766228 lpclm = 2.49779650178066e-7
+ pdiblc1 = 0.60630129375168 lpdiblc1 = -2.22569262949166e-7
+ pdiblc2 = -9.79659804609995e-05 lpdiblc2 = 3.10881001099169e-10
+ pdiblcb = -0.025
+ drout = 0.823688067692801 ldrout = 8.69813760605692e-8
+ pscbe1 = 800000000.0
+ pscbe2 = 7.5146551626052e-09 lpscbe2 = 8.89239691428671e-16
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.77191165332441 lbeta0 = 1.28254385565648e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -1.746561140738e-10 lagidl = 2.7282635504184e-16 pagidl = 9.4039548065783e-38
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.51916168720948 lkt1 = 5.27954896455041e-9
+ kt2 = -0.0724470689491601 lkt2 = 8.51455455724071e-9
+ at = -18539.604612764 lat = 0.0412132614604518 pat = 1.32348898008484e-23
+ ute = -2.133537872814 lute = 9.33843384158313e-7
+ ua1 = -1.02651999654268e-09 lua1 = 7.80820851034373e-16 wua1 = 3.94430452610506e-31
+ ub1 = 4.09283428091281e-19 lub1 = 7.01657725323038e-26
+ uc1 = 7.02451467413761e-11 luc1 = -2.2656620043097e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.69 pmos
* DC IV MOS Parameters
+ lmin = 2.5e-07 lmax = 5e-07 wmin = 1e-06 wmax = 1.26e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.006443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.948890704288003+0*(0.007356/sqrt(l*w*mult))} lvth0 = -3.14813566396651e-9
+ k1 = 0.43987873475056 lk1 = 3.41566092897283e-8
+ k2 = 0.00505947892961119 lk2 = -4.76964670712773e-09 pk2 = 1.57772181044202e-30
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 30780.1582495202 lvsat = 0.0198460709948983
+ ua = -7.20111477664003e-10 lua = -2.01569037735197e-16
+ ub = 1.1641954604768e-18 lub = 1.26449603631697e-25
+ uc = -4.30670652829792e-11 luc = 1.04933423200104e-17
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.00915178201416 lu0 = -8.78428769701665e-10
+ a0 = 1.44987763288 la0 = -1.55193100249753e-7
+ keta = -0.0561205618279248 lketa = 1.12302716530708e-8
+ a1 = 0.0
+ a2 = 1.06891451743248 la2 = -1.32665750201105e-7
+ ags = 2.17978636967648 lags = -4.27784020941055e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.18456167847128+0*(0.0/sqrt(l*w*mult))} lvoff = -5.78235162615357e-8
+ nfactor = {1.356397574+0*(0.1/sqrt(l*w*mult))} lnfactor = 4.05401698337989e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.49
+ etab = 4.850105e-05 letab = -2.70107735049e-11 petab = 9.24446373305873e-33
+ dsub = 0.0151130540728808 ldsub = 1.49138754216033e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.615591804575359 lpclm = 5.24672630688115e-9
+ pdiblc1 = -0.14347143930832 lpdiblc1 = 1.47322117633188e-07 ppdiblc1 = -5.04870979341448e-29
+ pdiblc2 = -0.00972230637784599 lpdiblc2 = 5.05893384406429e-09 wpdiblc2 = 8.27180612553028e-25 ppdiblc2 = -1.97215226305253e-31
+ pdiblcb = 0.1696704 lpdiblcb = -9.60383057952e-08 wpdiblcb = -5.29395592033938e-23 ppdiblcb = 1.26217744835362e-29
+ drout = 1.55317580771432 ldrout = -2.72902646626167e-7
+ pscbe1 = 800069244.261281 lpscbe1 = -0.034160825371373
+ pscbe2 = 9.42176599694321e-09 lpscbe2 = -5.16105533619634e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.77756825213281 lbeta0 = 1.2546377042271e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 6.493122281476e-10 lagidl = -1.33668538972981e-16
+ bgidl = 730034204.006401 lbgidl = 133.18438586389
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.504946199280001 lkt1 = -1.73349141960335e-9
+ kt2 = -0.0917821417920001 lkt2 = 1.80532807233817e-8
+ at = 63485.4642880001 lat = 0.000747178019086636
+ ute = -0.29451476672 lute = 2.65834030441113e-8
+ ua1 = 7.0578500184e-10 lua1 = -7.3791032257742e-17
+ ub1 = 6.6102183352e-19 lub1 = -5.40263489250896e-26
+ uc1 = 4.74348323563201e-11 luc1 = -1.14034251650022e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.24e-6
+ sbref = 1.24e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.70 pmos
* DC IV MOS Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 1e-06 wmax = 1.26e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.006443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.758071657257144+0*(0.007356/sqrt(l*w*mult))} lvth0 = -4.95816609303614e-8
+ k1 = -0.777750412353429 lk1 = 3.30452050687719e-7
+ k2 = 0.462511999162372 lk2 = -1.16085228075527e-07 wk2 = -2.11758236813575e-22
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 237786.933100285 lvsat = -0.0305265435837374
+ ua = 1.09572681037143e-10 lua = -4.03462721545216e-16
+ ub = 3.70232301220002e-19 lub = 3.19651010878927e-25
+ uc = -3.747113248118e-13 luc = 1.04670292537848e-19 wuc = -1.92592994438724e-34 puc = 2.29588740394978e-41
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0106202771988571 lu0 = -1.2357694509555e-9
+ a0 = 0.131411673999997 la0 = 1.65639769252188e-7
+ keta = -0.101820143345726 lketa = 2.23507164204494e-08 wketa = 2.64697796016969e-23 pketa = 1.26217744835362e-29
+ a1 = 0.0
+ a2 = 0.119936524349429 la2 = 9.82566566797385e-8
+ ags = -1.62902379023886 lags = 4.99044225752423e-7
+ b0 = 0.0
+ b1 = -5.21832167044571e-24 lb1 = 1.26981595864292e-30
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.220178493333428+0*(0.0/sqrt(l*w*mult))} lvoff = -4.91565917666102e-8
+ nfactor = {0.873008799999994+0*(0.1/sqrt(l*w*mult))} lnfactor = 5.230285558256e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 1.17996084013057 leta0 = -1.67893690915693e-7
+ etab = 0.0779204436747429 letab = -1.89762135479246e-08 wetab = 2.35746474577613e-23 petab = 1.62702561701834e-30
+ dsub = 1.515770617532 ldsub = -2.16028255960982e-07 wdsub = -1.6940658945086e-21
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.674530623428858 lpclm = -9.09532799529139e-9
+ pdiblc1 = 1.228866610524 lpdiblc1 = -1.86619878736909e-07 ppdiblc1 = 2.01948391736579e-28
+ pdiblc2 = 0.03274100563686 lpdiblc2 = -5.27400357497024e-9
+ pdiblcb = -0.596438571428571 lpdiblcb = 9.03851190942857e-8
+ drout = -0.975627884694001 ldrout = 3.42451386277088e-7
+ pscbe1 = 799752699.066854 lpscbe1 = 0.0428666491488912
+ pscbe2 = 8.76724844606286e-09 lpscbe2 = 1.07658438434153e-16
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 10.5332516765828 lbeta0 = -3.01760722716119e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 1956850179.27428 lbgidl = -165.346559925846
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.20003683742857 lkt1 = -7.59295257138061e-8
+ kt2 = 0.235996541485714 lkt2 = -6.17077285080508e-08 wkt2 = 5.29395592033938e-23 pkt2 = 1.26217744835362e-29
+ at = 84910.017942857 lat = -0.00446623001817895
+ ute = -0.108778416857143 lute = -1.86133088588166e-8
+ ua1 = 1.02665585028571e-09 lua1 = -1.51871102776825e-16
+ ub1 = 4.39e-19
+ uc1 = -3.41423648285715e-13 luc1 = 2.22353418646549e-19
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.71 pmos
* DC IV MOS Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 1e-06 wmax = 1.26e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.006443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {0.0887006526805187+0*(0.007356/sqrt(l*w*mult))} lvth0 = -1.96359479590336e-07 wvth0 = -1.00780724473305e-06 pvth0 = 1.74691292187539e-13
+ k1 = 3.75173699010685 lk1 = -4.5468023667994e-07 wk1 = -4.60324701042119e-06 pk1 = 7.9791763029239e-13
+ k2 = -0.736579800550957 lk2 = 9.17629463031819e-08 wk2 = 1.10786283713848e-06 pk2 = -1.92034728463909e-13
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -323162.505808177 lvsat = 0.0667073102577777 wvsat = 0.542257297594787 pvsat = -9.39937954504853e-8
+ ua = -1.31393747733486e-08 lua = 1.89308333230309e-15 wua = 1.57221619003511e-14 pua = -2.72524809948305e-21
+ ub = 1.03322383706342e-17 lub = -1.4071431971812e-24 wub = -1.23257039325945e-23 pub = 2.13651286826807e-30
+ uc = 1.91739534997083e-12 luc = -2.92638894255624e-19 wuc = -1.78688383262543e-18 puc = 3.09734869779627e-25
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = -0.0253214631398974 lu0 = 4.99429993588354e-09 wu0 = 3.98074765936302e-08 pu0 = -6.90014837778667e-15
+ a0 = -1.68631396147731 la0 = 4.80720695454553e-07 wa0 = 4.72212773875486e-06 pa0 = -8.1852417798029e-13
+ keta = 0.642009079699266 lketa = -1.06583153443723e-07 wketa = -5.0754522297849e-07 pketa = 8.79768738606455e-14
+ a1 = 0.0
+ a2 = 2.22133314433735 la2 = -2.65995230635728e-07 wa2 = -3.17932310752062e-06 pa2 = 5.51097508811409e-13
+ ags = 1.25
+ b0 = 0.0
+ b1 = 1.21760838977067e-23 lb1 = -1.74529551372948e-30
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {0.241123253568276+0*(0.0/sqrt(l*w*mult))} lvoff = -1.29117713971058e-07 wvoff = -1.08920521429769e-06 pvoff = 1.88800653435934e-13
+ nfactor = {-9.87283685517585+0*(0.1/sqrt(l*w*mult))} lnfactor = 2.38569195000247e-06 wnfactor = 1.3553173135453e-05 pnfactor = -2.34927992495316e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 2.75461061823134 leta0 = -4.40840334152124e-07 weta0 = -3.32646882694641e-06 peta0 = 5.76603453525237e-13
+ etab = 0.172175835684881 letab = -3.53142546881779e-08 wetab = -3.72130626979222e-07 petab = 6.45043786193245e-14
+ dsub = 0.43612777627507 ldsub = -2.88851251431879e-08 wdsub = -1.58885784466345e-07 pdsub = 2.75409441078276e-14
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -2.48628077310331 lpclm = 5.38793397856802e-07 wpclm = 4.10715258037321e-06 ppclm = -7.11925613976732e-13
+ pdiblc1 = -2.16557451097412 lpdiblc1 = 4.01765756381333e-07 wpdiblc1 = 3.09889307556994e-06 ppdiblc1 = -5.37155927933143e-13
+ pdiblc2 = -0.0421335406898698 lpdiblc2 = 7.70460053621247e-09 wpdiblc2 = 5.6113190420557e-08 ppdiblc2 = -9.72654820111851e-15
+ pdiblcb = 3.22192240415097 lpdiblcb = -5.71481935690721e-07 wpdiblcb = -3.8369659952901e-06 ppdiblcb = 6.65092011691596e-13
+ drout = 1.0
+ pscbe1 = 800000000.0
+ pscbe2 = 1.41961622561841e-08 lpscbe2 = -8.33378623584643e-16 wpscbe2 = -4.98576554589766e-15 ppscbe2 = 8.64222628194804e-22
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = -0.376966146498177 lbeta0 = 1.5893946143011e-06 wbeta0 = 1.73551820565636e-05 pbeta0 = -3.00831254732062e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 8.67672932376725e-09 lagidl = -1.48667310752317e-15 wagidl = -1.31156041904019e-14 pagidl = 2.27343259915589e-21
+ bgidl = 1017064548.30667 lbgidl = -2.44599822518103
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.295597738666668 lkt1 = -5.93651902149972e-8
+ kt2 = -0.12
+ at = -477168.708323278 lat = 0.0929633722353404 wat = 0.753758361715837 pat = -1.306549669031e-7
+ ute = -0.233981691333334 lute = 3.08917633233733e-9
+ ua1 = -1.45964257110642e-09 lua1 = 2.79098892990444e-16 wua1 = 1.90530345781488e-15 pua1 = -3.30261490770716e-22
+ ub1 = 7.73885347333333e-19 lub1 = -5.80483563360657e-26
+ uc1 = 3.8082395871078e-12 luc1 = -4.96940907250094e-19 wuc1 = -3.82172392294229e-17 puc1 = 6.62449981354972e-24
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.72 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.004443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.0053647+0*(0.005856/sqrt(l*w*mult))}
+ k1 = 0.49177002
+ k2 = -0.002473247
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 55237.817
+ ua = -1.3943119e-9
+ ub = 1.565972e-18
+ uc = -3.8916596e-11
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0072382252
+ a0 = 1.248405
+ keta = 0.0066402373
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.25185017
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.29956891+0*(0.0/sqrt(l*w*mult))}
+ nfactor = {1.7720538+0*(0.1/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.0017402344
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00056783834
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 799985290.0
+ pscbe2 = 1.0771971e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.0
+ alpha1 = 0.0
+ beta0 = 30.0
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.4670794e-10
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.54561
+ kt2 = -0.052484
+ at = 10000.0
+ ute = -1.2595
+ ua1 = -2.5605e-10
+ ub1 = 4.9434e-19
+ uc1 = 8.1951e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.73 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.004443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.0053647+0*(0.005856/sqrt(l*w*mult))}
+ k1 = 0.49177002
+ k2 = -0.002473247
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 55237.817
+ ua = -1.3943119e-9
+ ub = 1.565972e-18
+ uc = -3.8916596e-11
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0072382252
+ a0 = 1.248405
+ keta = 0.0066402373
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.25185017
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.29956891+0*(0.0/sqrt(l*w*mult))}
+ nfactor = {1.7720538+0*(0.1/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.0017402344
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00056783834
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 799985290.0
+ pscbe2 = 1.0771971e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.0
+ alpha1 = 0.0
+ beta0 = 30.0
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.4670794e-10
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.54561
+ kt2 = -0.052484
+ at = 10000.0
+ ute = -1.2595
+ ua1 = -2.5605e-10
+ ub1 = 4.9434e-19
+ uc1 = 8.1951e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.74 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.004443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.0074140810616+0*(0.005856/sqrt(l*w*mult))} lvth0 = 1.63813955161632e-8
+ k1 = 0.533711539863404 lk1 = -3.35252744501908e-7
+ k2 = -0.015204835164966 lk2 = 1.01767887479373e-07 wk2 = -3.30872245021211e-24
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 67709.0584957215 lvsat = -0.0996868485549274
+ ua = -1.96104979334726e-09 lua = 4.53012753893265e-15
+ ub = 1.85327925148432e-18 lub = -2.29654397096517e-24
+ uc = -2.32886427786375e-11 luc = -1.24919512346539e-16
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.00467602486377941 lu0 = 2.04805333111249e-8
+ a0 = 1.3219165622399 la0 = -5.87602763891561e-7
+ keta = 0.0100523898791525 lketa = -2.72744888727377e-8
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.199837851034395 lags = 4.15752045655891e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.318274014675695+0*(0.0/sqrt(l*w*mult))} lvoff = 1.49516223998211e-7
+ nfactor = {1.4620747314211+0*(0.1/sqrt(l*w*mult))} lnfactor = 2.47776746807634e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.0344627685079662 lpclm = 2.89382838858357e-07 wpclm = 3.30872245021211e-24 ppclm = -2.52435489670724e-29
+ pdiblc1 = 0.39
+ pdiblc2 = 9.85732448773808e-05 lpdiblc2 = 3.75099451691725e-9
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 799970624.466194 lpscbe1 = 0.117226568647311
+ pscbe2 = 1.20389481292726e-08 lpscbe2 = -1.01273764325455e-14
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.0
+ alpha1 = 0.0
+ beta0 = 30.0
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.35955228517575e-10 lagidl = 8.59500572955037e-17
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.629799548385 lkt1 = 6.72955516308661e-7
+ kt2 = -0.078183126699 lkt2 = 2.05421806009932e-7
+ at = -35193.10531325 lat = 0.361243766038403 wat = 1.38777878078145e-17
+ ute = -2.44701888775 lute = 9.49223985116982e-6
+ ua1 = -2.428076454925e-09 lua1 = 1.73617415991573e-14 pua1 = -1.50463276905253e-36
+ ub1 = 2.00166536148e-18 lub1 = -1.20485610902818e-23 pub1 = 5.60519385729927e-45
+ uc1 = 9.624331106095e-11 luc1 = -7.03799111305513e-16 wuc1 = 1.23259516440783e-32 puc1 = 9.4039548065783e-38
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.75 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.004443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.0087865031501+0*(0.005856/sqrt(l*w*mult))} lvth0 = 2.1861940794213e-8
+ k1 = 0.43831917185229 lk1 = 4.56812235868587e-8
+ k2 = 0.01332183338898 lk2 = -1.21487420705046e-8
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 32089.6541526299 lvsat = 0.0425534723457046
+ ua = -6.30371477103069e-10 lua = -7.83720747101323e-16
+ ub = 1.12874327553622e-18 lub = 5.96773074155464e-25
+ uc = -6.40771220126369e-11 luc = 3.79626717408019e-17
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0104860229284 lu0 = -2.72075274025099e-9
+ a0 = 1.2151813426064 la0 = -1.61372955390757e-7
+ keta = 0.0112322389301054 lketa = -3.19860249221718e-08 pketa = -1.26217744835362e-29
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.231933635768609 lags = 2.87582728836931e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.28016803107749+0*(0.0/sqrt(l*w*mult))} lvoff = -2.65384833187881e-9
+ nfactor = {2.3908807178428+0*(0.1/sqrt(l*w*mult))} lnfactor = -1.23126877212893e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.1592351855 leta0 = -3.16412877194199e-7
+ etab = -0.139268494014963 letab = 2.76612509352725e-7
+ dsub = 0.8590007 ldsub = -1.1940108573366e-6
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.275233282675524 lpclm = 1.2508608823632e-06 wpclm = 1.05879118406788e-22 ppclm = -8.07793566946316e-28
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0018580315657347 lpdiblc2 = -3.27511725517847e-9
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 799999960.06662 lpscbe1 = 7.96007225289941e-5
+ pscbe2 = 9.63319118340849e-09 lpscbe2 = -5.20375801862541e-16
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -3.038830824303e-12 lalpha0 = 1.21350786062605e-17
+ alpha1 = 2.9141211206745e-15 lalpha1 = -1.16370706077921e-20
+ beta0 = 56.910063 lbeta0 = -0.000107460977160294
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 6.68775207909697e-11 lagidl = 3.6180069251305e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.451622277389999 lkt1 = -3.85665506919708e-8
+ kt2 = -0.00801757949699999 lkt2 = -7.4772939922609e-8
+ at = 102918.248221 lat = -0.190281550261352
+ ute = 0.75230175845 lute = -3.28372885948521e-06 wute = 3.17637355220363e-22
+ ua1 = 3.98560513679e-09 lua1 = -8.2502568209387e-15
+ ub1 = -2.77182014511e-18 lub1 = 7.01357997563327e-24 wub1 = -1.46936793852786e-39 pub1 = -2.80259692864963e-45
+ uc1 = -2.21393444354e-10 luc1 = 5.64631814289713e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.76 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.004443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.006776922084+0*(0.005856/sqrt(l*w*mult))} lvth0 = 1.78561664910766e-8
+ k1 = 0.46881085865252 lk1 = -1.50990143961371e-8
+ k2 = 0.00448373627148801 lk2 = 5.46857276148265e-9
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 77900.2948653419 lvsat = -0.0487626185912911
+ ua = -1.30087102961762e-09 lua = 5.52811489908926e-16
+ ub = 1.65098192376424e-18 lub = -4.44225068426085e-25
+ uc = -4.1409249958814e-11 luc = -7.22205900322166e-18
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.00867459456899999 lu0 = 8.90036242818685e-10
+ a0 = 1.6312399809578 la0 = -9.9071844944486e-7
+ keta = 0.0279922647790546 lketa = -6.53944213278646e-08 wketa = 6.61744490042422e-24
+ a1 = 0.0
+ a2 = 0.8
+ ags = -0.393439099563341 lags = 1.53416196633805e-6
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.2886710916924+0*(0.0/sqrt(l*w*mult))} lvoff = 1.42956255081255e-8
+ nfactor = {1.4973376453944+0*(0.1/sqrt(l*w*mult))} lnfactor = 5.49864588819217e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = -0.0784703710000001 leta0 = 1.57414641388398e-07 weta0 = -1.24077091882954e-23 peta0 = -2.52435489670724e-29
+ etab = 0.00595669402992638 letab = -1.2870376534299e-08 wetab = 1.65436122510606e-24 petab = -5.52202633654708e-30
+ dsub = -0.0380014000000002 ldsub = 5.94017514673201e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.33332554131772 lpclm = 3.77974532621582e-8
+ pdiblc1 = 0.39770896841646 lpdiblc1 = -1.53665796853292e-8
+ pdiblc2 = 0.000215
+ pdiblcb = -0.423667599999999 lpdiblcb = 3.960116764488e-7
+ drout = 0.2110872461536 ldrout = 6.95501050926675e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 1.032799802395e-08 lpscbe2 = -1.90536067977383e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -9.32561383513941e-11 lalpha0 = 1.91968665957697e-16 walpha0 = -4.93038065763132e-32 palpha0 = -8.81620763116716e-38
+ alpha1 = -9.93396282422415e-11 lalpha1 = 1.98011627638891e-16 walpha1 = 1.17301170675335e-32 palpha1 = 4.12628363674874e-38
+ beta0 = -2.86171356345561 lbeta0 = 1.16843763911515e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 3.9577639605148e-10 lagidl = -2.93805933700986e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.428378914775259 lkt1 = -8.48984286397136e-8
+ kt2 = -0.02730481378342 lkt2 = -3.63269629045852e-8
+ at = -7927.86288261801 lat = 0.030672215153712
+ ute = -0.598656317552999 lute = -5.90812790181536e-7
+ ua1 = -6.67381794886596e-11 lua1 = -1.72566899554434e-16
+ ub1 = 1.01168299679436e-18 lub1 = -5.28220610244075e-25
+ uc1 = 7.61992951773119e-11 luc1 = -2.85711019421528e-17 wuc1 = -9.86076131526265e-32
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.77 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.004443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.021883259604+0*(0.005856/sqrt(l*w*mult))} lvth0 = 3.28618655905177e-8
+ k1 = 0.39884624356388 lk1 = 5.43994964267828e-8
+ k2 = 0.0243921037457624 lk2 = -1.43071651686781e-8
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -12824.776391484 lvsat = 0.041358042240822 pvsat = -2.64697796016969e-23
+ ua = -3.65131486012761e-10 lua = -3.76694156856437e-16
+ ub = 9.89933100099277e-19 lub = 2.12419847975622e-25
+ uc = -7.52043260124921e-11 luc = 2.63478742537868e-17
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0117406951944 lu0 = -2.1556380202149e-09 wu0 = 1.32348898008484e-23
+ a0 = 0.139135158719601 la0 = 4.91445970467591e-7
+ keta = -0.0422650138775481 lketa = 4.39480333832778e-09 wketa = -5.29395592033938e-23
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.991513061907201 lags = 1.58436356167227e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.24715506755244+0*(0.0/sqrt(l*w*mult))} lvoff = -2.69438188790142e-8
+ nfactor = {1.92532561224+0*(0.1/sqrt(l*w*mult))} lnfactor = 1.24727877808744e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = -0.32453716 leta0 = 4.0184213344008e-07 weta0 = 1.05879118406788e-22 peta0 = -2.01948391736579e-28
+ etab = -0.013900565275 letab = 6.85459370913796e-9
+ dsub = 0.79934936382752 ldsub = -2.37754818365701e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.11992164766228 lpclm = 2.49779650178066e-7
+ pdiblc1 = 0.60630129375168 lpdiblc1 = -2.22569262949166e-7
+ pdiblc2 = -9.79659804609995e-05 lpdiblc2 = 3.10881001099169e-10 ppdiblc2 = -1.97215226305253e-31
+ pdiblcb = -0.025
+ drout = 0.8236880676928 ldrout = 8.69813760605692e-8
+ pscbe1 = 800000000.0
+ pscbe2 = 7.51465516260521e-09 lpscbe2 = 8.89239691428677e-16
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.77191165332439 lbeta0 = 1.28254385565641e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -1.746561140738e-10 lagidl = 2.72826355041841e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.519161687209481 lkt1 = 5.27954896455041e-9
+ kt2 = -0.07244706894916 lkt2 = 8.51455455724071e-9
+ at = -18539.604612764 lat = 0.0412132614604517
+ ute = -2.133537872814 lute = 9.33843384158313e-7
+ ua1 = -1.02651999654268e-09 lua1 = 7.80820851034374e-16 pua1 = 1.88079096131566e-37
+ ub1 = 4.0928342809128e-19 lub1 = 7.01657725323045e-26
+ uc1 = 7.0245146741376e-11 luc1 = -2.2656620043097e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.78 pmos
* DC IV MOS Parameters
+ lmin = 2.5e-07 lmax = 5e-07 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.006443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.948890704288001+0*(0.007356/sqrt(l*w*mult))} lvth0 = -3.14813566396651e-9
+ k1 = 0.43987873475056 lk1 = 3.41566092897283e-8
+ k2 = 0.00505947892961119 lk2 = -4.76964670712773e-9
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 30780.15824952 lvsat = 0.0198460709948983
+ ua = -7.20111477664003e-10 lua = -2.01569037735197e-16
+ ub = 1.1641954604768e-18 lub = 1.26449603631696e-25
+ uc = -4.30670652829792e-11 luc = 1.04933423200104e-17
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.00915178201416002 lu0 = -8.78428769701665e-10
+ a0 = 1.44987763288 la0 = -1.55193100249753e-7
+ keta = -0.0561205618279248 lketa = 1.12302716530708e-8
+ a1 = 0.0
+ a2 = 1.06891451743248 la2 = -1.32665750201105e-7
+ ags = 2.17978636967648 lags = -4.27784020941055e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.18456167847128+0*(0.0/sqrt(l*w*mult))} lvoff = -5.78235162615357e-8
+ nfactor = {1.35639757400001+0*(0.1/sqrt(l*w*mult))} lnfactor = 4.05401698337989e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.49
+ etab = 4.850105e-05 letab = -2.70107735049e-11 wetab = -1.29246970711411e-26 petab = 9.24446373305873e-33
+ dsub = 0.0151130540728799 ldsub = 1.49138754216033e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.615591804575361 lpclm = 5.24672630688115e-9
+ pdiblc1 = -0.14347143930832 lpdiblc1 = 1.47322117633188e-7
+ pdiblc2 = -0.009722306377846 lpdiblc2 = 5.05893384406429e-09 ppdiblc2 = 1.57772181044202e-30
+ pdiblcb = 0.1696704 lpdiblcb = -9.60383057952e-08 wpdiblcb = -1.05879118406788e-22 ppdiblcb = 5.04870979341448e-29
+ drout = 1.55317580771432 ldrout = -2.72902646626167e-7
+ pscbe1 = 800069244.26128 lpscbe1 = -0.0341608253716004
+ pscbe2 = 9.42176599694321e-09 lpscbe2 = -5.16105533619603e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.77756825213281 lbeta0 = 1.2546377042271e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 6.493122281476e-10 lagidl = -1.33668538972981e-16
+ bgidl = 730034204.006401 lbgidl = 133.184385863891
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.50494619928 lkt1 = -1.73349141960335e-9
+ kt2 = -0.0917821417920001 lkt2 = 1.80532807233817e-8
+ at = 63485.464288 lat = 0.000747178019086692
+ ute = -0.29451476672 lute = 2.65834030441114e-8
+ ua1 = 7.0578500184e-10 lua1 = -7.3791032257742e-17
+ ub1 = 6.61021833520001e-19 lub1 = -5.402634892509e-26
+ uc1 = 4.74348323563201e-11 luc1 = -1.14034251650022e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.24e-6
+ sbref = 1.24e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.79 pmos
* DC IV MOS Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.006443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.75807165725714+0*(0.007356/sqrt(l*w*mult))} lvth0 = -4.95816609303614e-8
+ k1 = -0.777750412353427 lk1 = 3.30452050687719e-7
+ k2 = 0.462511999162371 lk2 = -1.16085228075527e-07 wk2 = -5.29395592033938e-23 pk2 = -2.52435489670724e-29
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 237786.933100285 lvsat = -0.0305265435837373
+ ua = 1.09572681037143e-10 lua = -4.03462721545216e-16
+ ub = 3.70232301220002e-19 lub = 3.19651010878929e-25
+ uc = -3.74711324811799e-13 luc = 1.04670292537848e-19 puc = 2.29588740394978e-41
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0106202771988571 lu0 = -1.2357694509555e-9
+ a0 = 0.131411673999999 la0 = 1.65639769252188e-7
+ keta = -0.101820143345726 lketa = 2.23507164204494e-08 pketa = -6.31088724176809e-30
+ a1 = 0.0
+ a2 = 0.119936524349429 la2 = 9.82566566797391e-8
+ ags = -1.62902379023885 lags = 4.99044225752423e-7
+ b0 = 0.0
+ b1 = -5.21832167044571e-24 lb1 = 1.26981595864292e-30
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.22017849333343+0*(0.0/sqrt(l*w*mult))} lvoff = -4.91565917666104e-8
+ nfactor = {0.873008800000008+0*(0.1/sqrt(l*w*mult))} lnfactor = 5.23028555825598e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 1.17996084013057 leta0 = -1.67893690915693e-7
+ etab = 0.0779204436747427 letab = -1.89762135479246e-08 wetab = -3.30872245021211e-24 petab = -4.95503256091948e-30
+ dsub = 1.515770617532 ldsub = -2.16028255960982e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.674530623428856 lpclm = -9.09532799529139e-9
+ pdiblc1 = 1.228866610524 lpdiblc1 = -1.86619878736909e-7
+ pdiblc2 = 0.0327410056368599 lpdiblc2 = -5.27400357497024e-9
+ pdiblcb = -0.596438571428571 lpdiblcb = 9.03851190942857e-08 ppdiblcb = -1.0097419586829e-28
+ drout = -0.975627884693997 ldrout = 3.42451386277088e-7
+ pscbe1 = 799752699.066856 lpscbe1 = 0.0428666491493459
+ pscbe2 = 8.76724844606284e-09 lpscbe2 = 1.07658438434153e-16
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 10.5332516765829 lbeta0 = -3.01760722716119e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 1956850179.27428 lbgidl = -165.346559925845
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.20003683742857 lkt1 = -7.59295257138064e-8
+ kt2 = 0.235996541485714 lkt2 = -6.17077285080507e-08 wkt2 = 5.29395592033938e-23
+ at = 84910.017942857 lat = -0.00446623001817897
+ ute = -0.108778416857143 lute = -1.86133088588166e-8
+ ua1 = 1.02665585028571e-09 lua1 = -1.51871102776825e-16
+ ub1 = 4.39e-19
+ uc1 = -3.41423648285712e-13 luc1 = 2.22353418646549e-19
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.80 pmos
* DC IV MOS Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.006443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.68809962941481+0*(0.007356/sqrt(l*w*mult))} lvth0 = 1.11627527707503e-07 wvth0 = 8.57374992354309e-07 pvth0 = -1.48615666424711e-13
+ k1 = -4.79593045011757 lk1 = 1.02695534207368e-06 wk1 = 4.36960021314835e-06 pk1 = -7.57417761746708e-13
+ k2 = 0.774294181522594 lk2 = -1.70128928001483e-07 wk2 = -4.78165340726173e-07 pk2 = 8.28842238307933e-14
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 201423.849894585 lvsat = -0.0242234394670275 wvsat = -0.00842313753061186 pvsat = 1.46004981328121e-9
+ ua = 8.19003938326279e-09 lua = -1.80411465877561e-15 wua = -6.66822424112128e-15 pua = 1.15585665350748e-21
+ ub = -5.11203448390804e-18 lub = 1.26993617087945e-24 wub = 3.88680103113297e-24 pub = -6.73730317134527e-31
+ uc = -1.84786167456466e-12 luc = 3.60023227863309e-19 wuc = 2.16566535987591e-18 puc = -3.7539210215017e-25
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0302110942004943 lu0 = -4.63160248838528e-09 wu0 = -1.84873923204987e-08 pu0 = 3.2045676100506e-15
+ a0 = 11.3490942475238 la0 = -1.77881089267728e-06 wa0 = -8.96169035245999e-06 pa0 = 1.55340148231471e-12
+ keta = 2.73604915463084 lketa = -4.69559871952213e-07 wketa = -2.70574745812533e-06 pketa = 4.69008852896528e-13
+ a1 = 0.0
+ a2 = -0.807337235419329 la2 = 2.58988435650536e-7
+ ags = -16.580389915694 lags = 3.09068412720657e-06 wags = 1.87173127369585e-05 pags = -3.2444215551989e-12
+ b0 = 0.0
+ b1 = 1.21760838977067e-23 lb1 = -1.74529551372948e-30
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.7617021702891+0*(0.0/sqrt(l*w*mult))} lvoff = 2.18048039349531e-07 wvoff = 1.01324515235828e-06 pvoff = -1.75633888219479e-13
+ nfactor = {38.5196597012058+0*(0.1/sqrt(l*w*mult))} lnfactor = -6.00256661808762e-06 wnfactor = -3.72464726631354e-05 pnfactor = 6.45622907848257e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 1.16073378506698 leta0 = -1.6456091164508e-07 weta0 = -1.65330905357142e-06 peta0 = 2.86581284727963e-13
+ etab = -1.2852994633915 letab = 2.17321598703125e-07 wetab = 1.15784269991888e-06 petab = -2.00698137918539e-13
+ dsub = 0.11768710587126 ldsub = 2.63127437832675e-08 wdsub = 1.75394825452823e-07 pdsub = -3.04025882543413e-14
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -3.04834640137308 lpclm = 6.36220729729829e-07 wpclm = 4.69717658953751e-06 ppclm = -8.14199195677253e-13
+ pdiblc1 = 0.786477026603333 lpdiblc1 = -1.09936953039269e-7
+ pdiblc2 = 0.01132071733706 lpdiblc2 = -1.5610536416595e-9
+ pdiblcb = -0.43322835123459 lpdiblcb = 6.20945859463013e-8
+ drout = 1.0
+ pscbe1 = -22426056.9391708 lpscbe1 = 142.557687857722 wpscbe1 = 863.33533834865 ppscbe1 = -0.000149648820878678
+ pscbe2 = -5.82203873378868e-09 lpscbe2 = 2.63653629961527e-15 wpscbe2 = 1.60281848013586e-14 ppscbe2 = -2.77829349709789e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 16.4098268772649 lbeta0 = -1.32039451485194e-06 wbeta0 = -2.66622983146096e-07 pbeta0 = 4.62158946525801e-14
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -2.23766860745942e-08 lagidl = 3.896063810798e-15 wagidl = 1.94824764073878e-14 pagidl = -3.37705349550379e-21
+ bgidl = 1017064548.30666 lbgidl = -2.44599822518103
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.295597738666672 lkt1 = -5.93651902149972e-8
+ kt2 = -0.12
+ at = 240872.694333334 lat = -0.0315004884183513
+ ute = -0.233981691333334 lute = 3.08917633233733e-9
+ ua1 = 3.55377781333335e-10 lua1 = -3.55131048607573e-17
+ ub1 = 7.73885347333335e-19 lub1 = -5.8048356336065e-26
+ uc1 = -3.25980697233334e-11 luc1 = 5.81365593600315e-18 wuc1 = -6.16297582203915e-33 puc1 = -2.93873587705572e-39
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.81 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 6.4e-07 wmax = 8.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.004443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.965665208194601+0*(0.005856/sqrt(l*w*mult))} wvth0 = -3.53223131778187e-8
+ k1 = 0.53696217035377 wk1 = -4.02093632784939e-8
+ k2 = 0.0032854709802425 wk2 = -5.12377440492052e-9
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 161274.634028667 wvsat = -0.0943454308640837
+ ua = -3.06755650285381e-09 wua = 1.48875633408128e-15
+ ub = 2.14389095287385e-18 wub = -5.14198880551676e-25
+ uc = 6.14166013797161e-11 wuc = -8.92706797696628e-17
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = -0.0033077195627891 wu0 = 9.38317209432245e-9
+ a0 = 1.2396907970452 wa0 = 7.75339410825026e-9
+ keta = 0.0039938051129965 wketa = 2.3546423962153e-9
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.31008900098943 wags = -5.18175456099637e-8
+ b0 = 7.3488582699e-08 wb0 = -6.53858932454902e-14
+ b1 = -7.7516677147e-09 wb1 = 6.89698588614615e-15
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.13114231410195+0*(0.0/sqrt(l*w*mult))} wvoff = -1.49856249972842e-7
+ nfactor = {0.738744457629098+0*(0.1/sqrt(l*w*mult))} wnfactor = 9.19378927561639e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.0017402344
+ pdiblc1 = 0.39
+ pdiblc2 = -0.00036344016320659 wpdiblc2 = 8.28597784255739e-10
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 834086075.39378 wpscbe1 = -30.3409078179893
+ pscbe2 = 1.50971808672986e-08 wpscbe2 = -3.84832174279197e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -3.448711e-10 walpha0 = 3.0684637123042e-16
+ alpha1 = -3.448711e-10 walpha1 = 3.0684637123042e-16
+ beta0 = 123.115197 wbeta0 = -8.28485202322134e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -3.39325340101386e-09 wagidl = 3.14965299146862e-15
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.61458422 wkt1 = 6.13692742460839e-8
+ kt2 = -0.052484
+ at = 10000.0
+ ute = -1.2595
+ ua1 = -2.5605e-10
+ ub1 = 4.9434e-19
+ uc1 = 8.1951e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.82 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 6.4e-07 wmax = 8.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.004443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.9656652081946+0*(0.005856/sqrt(l*w*mult))} wvth0 = -3.53223131778196e-8
+ k1 = 0.53696217035377 wk1 = -4.02093632784945e-8
+ k2 = 0.0032854709802425 wk2 = -5.12377440492052e-9
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 161274.634028667 wvsat = -0.0943454308640837
+ ua = -3.06755650285381e-09 wua = 1.48875633408128e-15
+ ub = 2.14389095287385e-18 wub = -5.14198880551675e-25
+ uc = 6.1416601379716e-11 wuc = -8.92706797696628e-17
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = -0.0033077195627891 wu0 = 9.38317209432245e-9
+ a0 = 1.2396907970452 wa0 = 7.75339410825026e-9
+ keta = 0.0039938051129965 wketa = 2.35464239621531e-9
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.31008900098943 wags = -5.18175456099636e-8
+ b0 = 7.34885826990001e-08 wb0 = -6.53858932454902e-14
+ b1 = -7.7516677147e-09 wb1 = 6.89698588614615e-15
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.13114231410195+0*(0.0/sqrt(l*w*mult))} wvoff = -1.49856249972842e-7
+ nfactor = {0.738744457629098+0*(0.1/sqrt(l*w*mult))} wnfactor = 9.19378927561638e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.0017402344
+ pdiblc1 = 0.39
+ pdiblc2 = -0.00036344016320659 wpdiblc2 = 8.28597784255739e-10
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 834086075.393781 wpscbe1 = -30.3409078179893
+ pscbe2 = 1.50971808672986e-08 wpscbe2 = -3.84832174279196e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -3.448711e-10 walpha0 = 3.0684637123042e-16
+ alpha1 = -3.448711e-10 walpha1 = 3.0684637123042e-16
+ beta0 = 123.115197 wbeta0 = -8.28485202322134e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -3.39325340101386e-09 wagidl = 3.14965299146862e-15
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.614584219999999 wkt1 = 6.13692742460839e-8
+ kt2 = -0.052484
+ at = 10000.0
+ ute = -1.2595
+ ua1 = -2.5605e-10
+ ub1 = 4.9434e-19
+ uc1 = 8.1951e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.83 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 6.4e-07 wmax = 8.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.004443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.72515996207783+0*(0.005856/sqrt(l*w*mult))} lvth0 = -1.92243972298452e-06 wvth0 = -2.5113340078368e-07 pvth0 = 1.72505096738126e-12
+ k1 = 0.667501357871833 lk1 = -1.04344384807726e-06 wk1 = -1.19038447012418e-07 pk1 = 6.3010751051556e-13
+ k2 = 0.0446385709964666 lk2 = -3.30549305777485e-07 wk2 = -5.32452038535666e-08 pk2 = 3.84650850626182e-13
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 256146.501807898 lvsat = -0.7583429058507 wvsat = -0.167660745374951 pvsat = 5.86034089461667e-7
+ ua = -5.3916837571497e-09 lua = 1.8577534698599e-14 wua = 3.0523798103483e-15 pua = -1.24985709505373e-20
+ ub = 5.90316992781693e-19 lub = 1.24182417710151e-23 wub = 1.12371081857504e-24 pub = -1.30923658385982e-29
+ uc = 1.14852851320696e-10 luc = -4.27134007230733e-16 wuc = -1.22910316871228e-16 puc = 2.68892989550151e-22
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = -0.0284101931192186 lu0 = 2.00652555772603e-07 wu0 = 2.94382043778722e-08 pu0 = -1.60306651643325e-13
+ a0 = 1.55649481432839 la0 = -2.53232158990239e-06 wa0 = -2.08714170085369e-07 pa0 = 1.7302984066363e-12
+ keta = 0.0303000374491662 lketa = -2.10274606569534e-07 wketa = -1.80151864937686e-08 pketa = 1.62822927319806e-13
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.075526637590849 lags = 1.87493625272369e-06 wags = 1.10604932533931e-07 pags = -1.29829776660176e-12
+ b0 = 4.65955853583017e-07 lb0 = -3.13712355011351e-12 wb0 = -4.14580586269831e-13 pb0 = 2.7912312091498e-18
+ b1 = -1.65368460393553e-08 lb1 = 7.02228997392437e-14 wb1 = 1.47135297761173e-14 pb1 = -6.24802773043741e-20
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {0.118207338180848+0*(0.0/sqrt(l*w*mult))} lvoff = -1.99313605087888e-06 wvoff = -3.88355879149557e-07 pvoff = 1.90640814888414e-12
+ nfactor = {-1.9804230014034+0*(0.1/sqrt(l*w*mult))} lnfactor = 2.17352245786479e-05 wnfactor = 3.06293550629829e-06 pnfactor = -1.71341722559656e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.21129242978291 lpclm = -9.6683595263376e-06 wpclm = -1.10840097078876e-06 ppclm = 8.85982359904266e-12
+ pdiblc1 = 0.39
+ pdiblc2 = -0.00385536529229361 lpdiblc2 = 2.79121378274862e-08 wpdiblc2 = 3.5179859727273e-09 ppdiblc2 = -2.14971888036609e-14
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 868115469.255025 lpscbe1 = -272.008447068059 wpscbe1 = -60.6313441210723 ppscbe1 = 0.000242121695538007
+ pscbe2 = 2.09454004135187e-08 lpscbe2 = -4.67467955311434e-14 wpscbe2 = -7.92444644958011e-15 ppscbe2 = 3.25818425115085e-20
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -6.15893687774676e-10 lalpha0 = 2.16637514971765e-15 walpha0 = 5.47986604726753e-16 palpha0 = -1.92751539173511e-21
+ alpha1 = -6.89167701418303e-10 lalpha1 = 2.75207910738777e-15 walpha1 = 6.13181586828864e-16 palpha1 = -2.44864091958123e-21
+ beta0 = 194.26704357092 lbeta0 = -0.000568740758965504 wbeta0 = -0.000146155320734286 pbeta0 = 5.06032654111637e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -7.13596854634974e-09 lagidl = 2.99167871943888e-14 wagidl = 6.47013745768275e-15 pagidl = -2.65417546621991e-20
+ bgidl = 2107368073.11315 lbgidl = -8851.56729880212 wbgidl = -985.272105581455 pbgidl = 0.00787561296188425
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.532375164970481 lkt1 = -6.57124763511551e-07 wkt1 = -8.66825852328784e-08 pkt1 = 1.18342855434385e-12
+ kt2 = -0.187620131271737 lkt2 = 1.08018877326737e-06 wkt2 = 9.73707212099572e-08 pkt2 = -7.78317085934957e-13
+ at = -9258.91033287105 lat = 0.153942979802331 wat = -0.0230747476970713 pat = 1.84444257607413e-7
+ ute = -3.4587347911921 lute = 1.75792270273579e-05 wute = 9.00166333703561e-07 pute = -7.19533376151336e-12
+ ua1 = -7.74708200901268e-09 lua1 = 5.98783508168574e-14 wua1 = 4.73254370350619e-15 pua1 = -3.78288214218968e-20
+ ub1 = 6.95549342879971e-18 lub1 = -5.1646183226255e-23 wub1 = -4.40762988303878e-24 pub1 = 3.52316754340295e-29
+ uc1 = 2.18816134008649e-10 luc1 = -1.68356511474062e-15 wuc1 = -1.09058213149696e-16 puc1 = 8.71739159381564e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.84 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 6.4e-07 wmax = 8.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.004443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.48369657877072+0*(0.005856/sqrt(l*w*mult))} lvth0 = 1.10665337284664e-06 wvth0 = 4.22547535484859e-07 pvth0 = -9.65184715295479e-13
+ k1 = 0.310784755338068 lk1 = 3.81046116051721e-07 wk1 = 1.1347275232508e-07 pk1 = -2.98388297224449e-13
+ k2 = -0.0809058222230736 lk2 = 1.70791890353048e-07 wk2 = 8.38383216051109e-08 pk2 = -1.62770000761923e-13
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 6328.02789852174 lvsat = 0.23926669911362 wvsat = 0.022921206018908 pvsat = -1.75024059153584e-7
+ ua = 9.28935636043634e-10 lua = -6.66283490777689e-15 wua = -1.3873813413268e-15 pua = 5.23089596737064e-21
+ ub = 5.29866001719286e-18 lub = -6.38376334540092e-24 wub = -3.71015089553841e-24 pub = 6.21087783111622e-30
+ uc = -1.28738524394411e-11 luc = 8.29218925093662e-17 wuc = -4.55577097172483e-17 puc = -4.00021159969081e-23
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0423301789367373 lu0 = -8.1837660092584e-08 wu0 = -2.83330894240013e-08 pu0 = 7.0393651204861e-14
+ a0 = 0.805977799876988 la0 = 4.6474652355295e-07 wa0 = 3.64085660355861e-07 pa0 = -5.57084922658227e-13
+ keta = -0.0415269255683224 lketa = 7.65547342727979e-08 wketa = 4.6942055090993e-08 pketa = -9.65732938758026e-14
+ a1 = 0.0
+ a2 = 0.8
+ ags = 1.38197925172107 lags = -3.34217061648187e-06 wags = -1.0232441164379e-06 pags = 3.22954472692131e-12
+ b0 = -7.0518677536023e-07 lb0 = 1.53964481346546e-12 wb0 = 6.27434432919917e-13 pb0 = -1.36988696355135e-18
+ b1 = 3.32697706660904e-09 lb1 = -9.10005989508186e-15 wb1 = -2.96015189459428e-15 pb1 = 8.09670731118191e-21
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.564367221686601+0*(0.0/sqrt(l*w*mult))} lvoff = 7.32614876873084e-07 wvoff = 2.5286401309077e-07 pvoff = -6.54199613155058e-13
+ nfactor = {6.67145586754464+0*(0.1/sqrt(l*w*mult))} lnfactor = -1.28146520801193e-05 wnfactor = -3.80860835096105e-06 pnfactor = 1.03062249478946e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.1592351855 leta0 = -3.16412877194199e-7
+ etab = -0.1392684888935 letab = 2.76612488900993e-07 wetab = -4.55678155815718e-15 petab = 1.81967689549841e-20
+ dsub = 0.859000699999999 ldsub = -1.1940108573366e-6
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -2.94416912670563 lpclm = 6.92580301472722e-06 wpclm = 2.3746648495262e-06 ppclm = -5.04923549772225e-12
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00629790356823405 lpdiblc2 = -1.26332965374756e-08 wpdiblc2 = -3.95034148322218e-09 ppdiblc2 = 8.3263670226255e-15
+ pdiblcb = 0.462444668731799 lpdiblcb = -2.74519891854411e-06 wpdiblcb = -6.11648531935703e-07 ppdiblcb = 2.44251932522306e-12
+ drout = 0.56
+ pscbe1 = 799999822.347933 lpscbe1 = 0.000354120616975706 wpscbe1 = 0.000122534127513063 ppscbe1 = -2.44251931180717e-10
+ pscbe2 = 9.64315525817299e-09 lpscbe2 = -1.61311046698578e-15 wpscbe2 = -8.86545780193426e-18 ppscbe2 = 9.72252144963023e-22
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -1.47298006479066e-10 lalpha0 = 2.95114208964001e-16 walpha0 = 1.28353476317255e-16 palpha0 = -2.51778473998583e-22
+ alpha1 = 1.09856605183185e-14 lalpha1 = -4.43325141949713e-20 walpha1 = -7.18158922104643e-21 palpha1 = 2.90905159072328e-26
+ beta0 = 100.526597136953 lbeta0 = -0.00019440347208378 wbeta0 = -3.88074710393879e-05 pbeta0 = 7.73564067067115e-11
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 8.18678047687567e-10 lagidl = -1.84880532615097e-15 wagidl = -6.68908654762138e-16 pagidl = 1.96686946237936e-21
+ bgidl = -1214736146.2263 lbgidl = 4414.71772024643 wbgidl = 1970.54421116291 pbgidl = -0.00392796065679104
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.990108369035007 lkt1 = 1.17075863414108e-06 wkt1 = 4.7911379984963e-07 pkt1 = -1.07598765046876e-12
+ kt2 = 0.169707816943784 lkt2 = -3.46742500803708e-07 wkt2 = -1.58129785225095e-07 pkt2 = 2.41982795431383e-13
+ at = 162669.829780976 lat = -0.532626591386421 wat = -0.0531635036306529 pat = 3.0459883004971e-7
+ ute = 2.53384282221434 lute = -6.35116087420737e-06 wute = -1.58511226546402e-06 pute = 2.72922370912933e-12
+ ua1 = 1.51200806020696e-08 lua1 = -3.14379585901566e-14 wua1 = -9.90681269632386e-15 pua1 = 2.06310767850878e-20
+ ub1 = -1.34715955358992e-17 lub1 = 2.9926087365858e-23 wub1 = 9.52004169570669e-24 pub1 = -2.03862247328948e-29
+ uc1 = -5.20614354072123e-10 luc1 = 1.26923075167087e-15 wuc1 = 2.66229470498604e-16 puc1 = -6.26911408663171e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.85 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 6.4e-07 wmax = 8.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.004443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.859423135614458+0*(0.005856/sqrt(l*w*mult))} lvth0 = -1.37734603787577e-07 wvth0 = -1.3110688215174e-07 pvth0 = 1.38435674247424e-13
+ k1 = 0.657368028317915 lk1 = -3.09811492143383e-07 wk1 = -1.67767270963862e-07 pk1 = 2.62218128318286e-13
+ k2 = -0.0455948556104336 lk2 = 1.00405198787341e-07 wk2 = 4.4557036513923e-08 pk2 = -8.44691225008245e-14
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 762849.569148904 lvsat = -1.26873643687933 wvsat = -0.60942827418946 pvsat = 1.085462189026e-6
+ ua = -4.96352633601228e-09 lua = 5.0828334546771e-15 wua = 3.25881899015326e-15 pua = -4.03055170898115e-21
+ ub = 3.13693157806079e-18 lub = -2.07470790199829e-24 wub = -1.32211211450305e-24 pub = 1.45070938340477e-30
+ uc = 1.86582307318966e-10 luc = -3.14661650071138e-16 wuc = -2.02853709753758e-16 puc = 2.73541978123868e-22
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = -0.0099876454102004 lu0 = 2.24494472554921e-08 wu0 = 1.66045824560217e-08 pu0 = -1.91823177851203e-14
+ a0 = 3.45437665409091 la0 = -4.81440755170812e-06 wa0 = -1.62212163445413e-06 pa0 = 3.40209755396374e-12
+ keta = 0.163032746319274 lketa = -3.3120183296828e-07 wketa = -1.20151215134654e-07 pketa = 2.36500071209249e-13
+ a1 = 0.0
+ a2 = -0.570294274927202 la2 = 2.73145964939484e-06 wa2 = 1.21920864282113e-06 pa2 = -2.43029491766379e-12
+ ags = -4.12625971097633 lags = 7.63761142094344e-06 wags = 3.32124802300394e-06 pags = -5.4304965453294e-12
+ b0 = 5.57355890638085e-07 lb0 = -9.77029459290286e-13 wb0 = -4.95903056319289e-13 pb0 = 8.6930434057375e-19
+ b1 = -9.72774657807711e-09 lb1 = 1.69224168253695e-14 wb1 = 8.6551866414208e-15 pb1 = -1.50565883755213e-20
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0691986110760774+0*(0.0/sqrt(l*w*mult))} lvoff = -2.54423531064076e-07 wvoff = -1.95273927743024e-07 pvoff = 2.39090773550695e-13
+ nfactor = {7.84014345782272+0*(0.1/sqrt(l*w*mult))} lnfactor = -1.5144241463949e-05 wnfactor = -5.64346199772277e-06 pnfactor = 1.39637084464233e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 1.32608126080038 leta0 = -2.64233149924131e-06 weta0 = -1.24968885889166e-06 peta0 = 2.49105229060539e-12
+ etab = -0.535309554809244 letab = 1.06605619515135e-06 wetab = 4.81587423027911e-07 petab = -9.59966501530046e-13
+ dsub = -1.0657221061954 ldsub = 2.64261225171933e-06 wdsub = 9.1440648211585e-07 pdsub = -1.82272118824784e-12
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.73893377609808 lpclm = -2.40920395934172e-06 wpclm = -1.25062896315159e-06 ppclm = 2.17720042025328e-12
+ pdiblc1 = 0.426036787903175 lpdiblc1 = -7.18334987253389e-08 wpdiblc1 = -2.52044564313128e-08 ppdiblc1 = 5.02410007738801e-14
+ pdiblc2 = 0.00044351946819426 lpdiblc2 = -9.6353024427052e-10 wpdiblc2 = -2.03323414373991e-10 ppdiblc2 = 8.5729351930379e-16
+ pdiblcb = -2.4837040749272 lpdiblcb = 3.12747132584364e-06 wpdiblcb = 1.83290138528197e-06 ppdiblcb = -2.43029491766379e-12
+ drout = 0.132697301170835 ldrout = 8.51758707078729e-07 wdrout = 6.97468421068433e-08 pdrout = -1.39029030751571e-13
+ pscbe1 = 795876407.695818 lpscbe1 = 8.21971323643265 wpscbe1 = 3.66893408862597 ppscbe1 = -7.31342573835267e-6
+ pscbe2 = 1.13026784410869e-08 lpscbe2 = -4.92110108936893e-15 wpscbe2 = -8.67214298640282e-16 ppscbe2 = 2.68323150666203e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -9.78343046749665e-11 lalpha0 = 1.96516332537222e-16 walpha0 = 4.0733877767013e-18 palpha0 = -4.04625086733295e-24
+ alpha1 = -9.93562343796287e-11 lalpha1 = 1.98028123146192e-16 walpha1 = 1.47751812125238e-20 palpha1 = -1.4676748955295e-26
+ beta0 = -6.20685847615589 lbeta0 = 1.83523808611436e-05 wbeta0 = 2.97631659394476e-06 pbeta0 = -5.93280496674065e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.49936455062403e-09 lagidl = -3.20564359854133e-15 wagidl = -9.81908952543322e-16 pagidl = 2.59078484995791e-21
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.308869546253552 lkt1 = -1.87180598384462e-07 wkt1 = -1.06332528469114e-07 pkt1 = 9.10047627294653e-14
+ kt2 = 0.0692276212061779 lkt2 = -1.464515083925e-07 wkt2 = -8.58889810790018e-08 pkt2 = 9.79824553764174e-14
+ at = -60385.6255734575 lat = -0.0880016761211245 wat = 0.0466738851836254 pat = 1.05589169105434e-7
+ ute = 3.35565372383641 lute = -7.98930777322491e-06 wute = -3.5183165157079e-06 pute = 6.58275320290197e-12
+ ua1 = 3.20082681823455e-09 lua1 = -7.67885709119445e-15 wua1 = -2.90729046971724e-15 pua1 = 6.67866314894821e-21
+ ub1 = -7.15013116341382e-19 lub1 = 4.49790687882139e-24 wub1 = 1.53631439843284e-24 pub1 = -4.47195772960159e-30
+ uc1 = 1.29507157777217e-11 luc1 = 2.0565522246652e-16 wuc1 = 5.62749301818661e-17 puc1 = -2.08401045177286e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.86 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 6.4e-07 wmax = 8.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.004443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.02429016494824+0*(0.005856/sqrt(l*w*mult))} lvth0 = 2.6034081396777e-08 wvth0 = 2.14152525617169e-09 pvth0 = 6.07496772966427e-15
+ k1 = 0.277808267571465 lk1 = 6.72196414769748e-08 wk1 = 1.07692595043038e-07 pk1 = -1.14066240612767e-14
+ k2 = 0.0902011196598536 lk2 = -3.44861036956955e-08 wk2 = -5.85530585992385e-08 pk2 = 1.79540531586932e-14
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -1028975.22170011 lvsat = 0.511151217213039 wvsat = 0.904111932739872 pvsat = -4.17994813044765e-7
+ ua = -8.66142550562498e-10 lua = 1.01274644000598e-15 wua = 4.45770686796826e-16 pua = -1.23624393342168e-21
+ ub = 2.1933894081532e-18 lub = -1.13745161002662e-24 wub = -1.07076586313177e-24 pub = 1.20103760076012e-30
+ uc = -2.07502846058195e-10 luc = 7.67981080142249e-17 wuc = 1.17711576282208e-16 puc = -4.48877019765265e-23
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.011010498421116 lu0 = 1.59119305837996e-09 wu0 = 6.49686883494607e-10 pu0 = -3.33371372689737e-15
+ a0 = -3.99208702022471 la0 = 2.58244778160921e-06 wa0 = 3.67572271018271e-06 pa0 = -1.86045255164913e-12
+ keta = -0.223389161120479 lketa = 5.26457317241094e-08 wketa = 1.61153797241049e-07 pketa = -4.29308871740078e-14
+ a1 = 0.0
+ a2 = 3.5405885498544 la2 = -1.35203647400807e-06 wa2 = -2.43841728564227e-06 pa2 = 1.20296390686419e-12
+ ags = 4.15204655216979 lags = -5.85544765877597e-07 wags = -2.81206002079992e-06 pags = 6.6195140028663e-13
+ b0 = -7.63776618893518e-07 lb0 = 3.35301665462817e-13 wb0 = 6.7956428920288e-13 pb0 = -2.98332041492551e-19
+ b1 = 7.07121378167302e-08 lb1 = -6.29815770595996e-14 wb1 = -6.29155730677607e-14 pb1 = 5.60373669324776e-20
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.502899797474587+0*(0.0/sqrt(l*w*mult))} lvoff = 1.76388338030647e-07 wvoff = 2.27546878639337e-07 pvoff = -1.80913200619547e-13
+ nfactor = {-16.2897037903437+0*(0.1/sqrt(l*w*mult))} lnfactor = 8.82485274185011e-06 wnfactor = 1.62066803337195e-05 pnfactor = -7.74086823680687e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = -3.13364042360076 leta0 = 1.78767951929836e-06 weta0 = 2.49937771778332e-06 peta0 = -1.23303800453579e-12
+ etab = 1.06863191191749 letab = -5.27199813524051e-07 wetab = -9.63174827828696e-07 petab = 4.75170743211353e-13
+ dsub = 2.78751565154149 ldsub = -1.18495523607552e-06 wdsub = -1.76895544679646e-06 pdsub = 8.42764183494051e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -1.96633750457257 lpclm = 1.27138280405711e-06 wpclm = 1.85623280787957e-06 ppclm = -9.08963437659276e-13
+ pdiblc1 = 0.689231955458777 lpdiblc1 = -3.33275260074686e-07 wpdiblc1 = -7.37869093947287e-08 ppdiblc1 = 9.84997974356532e-14
+ pdiblc2 = -0.000195366777709762 lpdiblc2 = -3.2890025853671e-10 wpdiblc2 = 8.66615996258679e-11 ppdiblc2 = 5.69240385467198e-16
+ pdiblcb = 0.6647422 wpdiblcb = -6.1369274246084e-7
+ drout = 0.420328173142241 ldrout = 5.66044031976397e-07 wdrout = 3.58886319969184e-07 pdrout = -4.26242261412392e-13
+ pscbe1 = 808247184.608363 lpscbe1 = -4.06864956032086 wpscbe1 = -7.33786817725104 ppscbe1 = 3.62004921082874e-6
+ pscbe2 = -2.48817233168534e-08 lpscbe2 = 3.102224018406e-14 wpscbe2 = 2.88244250603462e-14 ppscbe2 = -2.68106021509148e-20
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 15.5543404033212 lbeta0 = -3.26384491139844e-06 wbeta0 = -6.03461307736544e-06 pbeta0 = 3.01809389109928e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -3.97571285711779e-09 lagidl = 2.23295884351012e-15 wagidl = 3.3819605888808e-15 pagidl = -1.74401259258124e-21
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.489498227233902 lkt1 = -7.75526567680261e-09 wkt1 = -2.63928321382829e-08 pkt1 = 1.15976246555895e-14
+ kt2 = -0.170374632876666 lkt2 = 9.15545154736435e-08 wkt2 = 8.71302861694994e-08 pkt2 = -7.38841575136742e-14
+ at = -357041.480976851 lat = 0.206677857973572 wat = 0.301179404180311 pat = -1.47220834123696e-7
+ ute = -8.56891076383874 lute = 3.85581526583335e-06 wute = 5.72582283388071e-06 pute = -2.59980169033969e-12
+ ua1 = -1.03770323445347e-08 lua1 = 5.80854637383246e-15 wua1 = 8.31954542762961e-15 pua1 = -4.47337956765052e-21
+ ub1 = 6.77754494824054e-18 lub1 = -2.94473576393429e-24 wub1 = -5.66611101511295e-24 pub1 = 2.68248512583916e-30
+ uc1 = 4.13043360831461e-10 luc1 = -1.91772005385871e-16 wuc1 = -3.05002037160583e-16 puc1 = 1.50469095008728e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.87 pmos
* DC IV MOS Parameters
+ lmin = 2.5e-07 lmax = 5e-07 wmin = 6.4e-07 wmax = 8.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.006443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.980951512537821+0*(0.007356/sqrt(l*w*mult))} lvth0 = 4.65347729392831e-09 wvth0 = 2.85258540659735e-08 pvth0 = -6.94142427670586e-15
+ k1 = 0.252308782950744 lk1 = 7.97995062207916e-08 wk1 = 1.66888901568262e-07 pk1 = -4.06104115298177e-14
+ k2 = 0.0542080779936456 lk2 = -1.67293685061717e-08 wk2 = -4.37295826581519e-08 pk2 = 1.06410691848694e-14
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -95269.655412271 lvsat = 0.0505187805517312 wvsat = 0.112151838517032 pvsat = -2.72908040810576e-8
+ ua = 3.84897972353431e-09 lua = -1.31340255245239e-15 wua = -4.06531325735483e-15 pua = 9.89245197418209e-22
+ ub = -1.86044745912135e-18 lub = 8.62460162400871e-25 wub = 2.69115244549768e-24 pub = -6.54859653782514e-31
+ uc = -1.02337679370456e-10 luc = 2.49161350108288e-17 wuc = 5.27355665735425e-17 puc = -1.28325672988727e-23
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0226981710655859 lu0 = -4.17477998869755e-09 wu0 = -1.20527939966716e-08 pu0 = 2.93290278556207e-15
+ a0 = 1.66152932818236 la0 = -2.06696000481239e-07 wa0 = -1.8831544501205e-07 pa0 = 4.58243037583423e-14
+ keta = -0.22053854649493 lketa = 5.12394152059706e-08 wketa = 1.46289619397188e-07 pketa = -3.55978234048729e-14
+ a1 = 0.0
+ a2 = 1.06891451743248 la2 = -1.32665750201105e-7
+ ags = 5.44070696557385 lags = -1.22128991690553e-06 wags = -2.90137866501904e-06 pags = 7.06015681588403e-13
+ b0 = -1.65993456595493e-07 lb0 = 4.03925157410342e-14 wb0 = 1.47691383256879e-13 pb0 = -3.59389258189624e-20
+ b1 = -1.12386369653478e-07 lb1 = 2.7347874418738e-14 wb1 = 9.99948957854986e-14 pb1 = -2.43325579506517e-20
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {0.124092574886034+0*(0.0/sqrt(l*w*mult))} lvoff = -1.32930824964998e-07 wvoff = -2.74622714421495e-07 pvoff = 6.68261420818977e-14
+ nfactor = {0.21223232851807+0*(0.1/sqrt(l*w*mult))} lnfactor = 6.83820580843069e-07 wnfactor = 1.01801210267863e-06 pnfactor = -2.47721029041613e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.49
+ etab = 4.850105e-05 letab = -2.70107735049e-11 wetab = -6.46234853557053e-27 petab = -3.08148791101958e-33
+ dsub = 0.14966330342655 ldsub = 1.16397565638811e-07 wdsub = -1.19715034870482e-07 pdsub = 2.91312171553135e-14
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.585080749510564 lpclm = 1.26712254242382e-08 wpclm = 2.71469732576727e-08 ppclm = -6.60589017857557e-15
+ pdiblc1 = -0.422644040669374 lpdiblc1 = 2.15255420103184e-07 wpdiblc1 = 2.48391644514707e-07 ppdiblc1 = -6.04431259929198e-14
+ pdiblc2 = -0.0124736374744419 lpdiblc2 = 5.72843725044776e-09 wpdiblc2 = 2.44797538281369e-09 ppdiblc2 = -5.95685433703119e-16
+ pdiblcb = 1.5307745498544 lpdiblcb = -4.2724666741247e-07 wpdiblcb = -1.21103180072058e-06 ppdiblcb = 2.94690056323745e-13
+ drout = 2.67345537674649 ldrout = -5.45509236395318e-07 wdrout = -9.96760008365738e-07 pdrout = 2.42549586915702e-13
+ pscbe1 = 800069244.26128 lpscbe1 = -0.0341608253711456
+ pscbe2 = 6.60243097022716e-08 lpscbe2 = -1.38251603335292e-14 wpscbe2 = -5.0361671761975e-14 ppscbe2 = 1.22549084832155e-20
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.59329040294026 lbeta0 = 1.70305573689528e-07 wbeta0 = 1.63959778951856e-07 pbeta0 = -3.98976446905875e-14
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 9.89019256021353e-10 lagidl = -2.16332167721724e-16 wagidl = -3.02251678335855e-16 pagidl = 7.35493189028902e-23
+ bgidl = 730034204.006402 lbgidl = 133.184385863891
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.498549009775686 lkt1 = -3.29017071920441e-09 wkt1 = -5.6918494633865e-09 pkt1 = 1.38504326472157e-15
+ kt2 = 0.0471321477421401 lkt2 = -1.57498446632769e-08 wkt2 = -1.23597905581543e-07 pkt2 = 3.00760671484015e-14
+ at = 57360.4956136553 lat = 0.0022376156463644 wat = 0.00544964310324264 pat = -1.32610525345685e-9
+ ute = -1.30588320526931 lute = 2.72687776143824e-07 wute = 8.9985717952543e-07 pute = -2.18969446351359e-13
+ ua1 = 2.36483485009753e-09 lua1 = -4.77500904233033e-16 wua1 = -1.47612666189832e-15 pua1 = 3.59197709653013e-22
+ ub1 = 1.16823729496324e-18 lub1 = -1.77451144881766e-25 wub1 = -4.51291000538526e-25 pub1 = 1.09816249489044e-31
+ uc1 = 4.743483235632e-11 luc1 = -1.14034251650022e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.24e-6
+ sbref = 1.24e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.88 pmos
* DC IV MOS Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 6.4e-07 wmax = 8.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.006443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.708437786079259+0*(0.007356/sqrt(l*w*mult))} lvth0 = -6.16594678750467e-08 wvth0 = -4.41613497363315e-08 pvth0 = 1.07461345221392e-14
+ k1 = -2.02711795768269 lk1 = 6.34470650433051e-07 wk1 = 1.11161502838986e-06 pk1 = -2.70498177778332e-13
+ k2 = 0.545014304567405 lk2 = -1.36161174068177e-07 wk2 = -7.34057827161471e-08 pk2 = 1.78624163545817e-14
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 738412.672293368 lvsat = -0.152347809707504 wvsat = -0.445427846566279 pvsat = 1.08389521327745e-7
+ ua = 5.86452439728656e-09 lua = -1.80386116227392e-15 wua = -5.12042340090954e-15 pua = 1.24599358953053e-21
+ ub = 1.32705326660253e-18 lub = 8.68201108046759e-26 wub = -8.51323990745568e-25 pub = 2.07159477260045e-31
+ uc = -1.68800651054782e-12 luc = 4.2424491644448e-19 wuc = 1.16849414780618e-18 puc = -2.8433902893886e-25
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0375241069894086 lu0 = -7.78249358452872e-09 wu0 = -2.39374727062708e-08 pu0 = 5.82489673339853e-15
+ a0 = 1.95638728836938 la0 = -2.78446146797227e-07 wa0 = -1.62375781807536e-06 pa0 = 3.95121979934823e-13
+ keta = 0.182152680668966 lketa = -4.67506626296377e-08 wketa = -2.52662605179045e-07 pketa = 6.14824130190584e-14
+ a1 = 0.0
+ a2 = -0.0353204792273516 la2 = 1.36036585416105e-07 wa2 = 1.38138707927813e-07 pa2 = -3.36143969097381e-14
+ ags = -1.62902379023885 lags = 4.99044225752423e-7
+ b0 = -4.26994762369998e-09 lb0 = 1.0390405148559e-15 wb0 = 3.79915259259559e-15 pb0 = -9.24478193577026e-22
+ b1 = 6.44215537882842e-10 lb1 = -1.56762120557335e-16 wb1 = -5.73185749950068e-16 pb1 = 1.3947787402135e-22
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {0.412683937009636+0*(0.0/sqrt(l*w*mult))} lvoff = -2.03156069841431e-07 wvoff = -5.63084411070787e-07 pvoff = 1.37019834421143e-13
+ nfactor = {23.1890864511252+0*(0.1/sqrt(l*w*mult))} lnfactor = -4.90732114764391e-06 wnfactor = -1.9855556024683e-05 pnfactor = 4.83161129193432e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.430993751557764 leta0 = 1.43584624834372e-08 weta0 = 6.66387625114366e-07 peta0 = -1.62157431920079e-13
+ etab = -0.497100985801246 letab = 1.20948351057903e-07 wetab = 5.11620831709111e-07 petab = -1.24496789946432e-13
+ dsub = 1.44415360420511 ldsub = -1.98601115172043e-07 wdsub = 6.37206789948942e-08 pdsub = -1.55056625852597e-14
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.708064400894729 lpclm = -1.72553703362815e-08 wpclm = -2.9836416936794e-08 ppclm = 7.26033402456562e-15
+ pdiblc1 = 1.37328460825487 lpdiblc1 = -2.21762265468745e-07 wpdiblc1 = -1.28494787020665e-07 ppdiblc1 = 3.12676644840345e-14
+ pdiblc2 = 0.0418517851956429 lpdiblc2 = -7.49100245124536e-09 wpdiblc2 = -8.10624504834657e-09 ppdiblc2 = 1.97255745757456e-15
+ pdiblcb = 0.0440041723303621 lpdiblcb = -6.54589372865257e-08 wpdiblcb = -5.6982893580611e-07 ppdiblcb = 1.38661033581187e-13
+ drout = -0.975627884693997 ldrout = 3.42451386277089e-7
+ pscbe1 = 799752699.066856 lpscbe1 = 0.0428666491488912
+ pscbe2 = -6.28682802277113e-08 lpscbe2 = 1.7539304714853e-14 wpscbe2 = 6.3737152880367e-14 ppscbe2 = -1.55096713076027e-20
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 6.97931790606873 lbeta0 = 5.63046413133249e-07 wbeta0 = 3.16208485163153e-06 pbeta0 = -7.69455403626315e-13
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 3.86620788894034e-08 lagidl = -9.38361915278965e-15 wagidl = -3.43103089076314e-14 pagidl = 8.3490019489652e-21
+ bgidl = 1931628452.65062 lbgidl = -159.209155412696 wbgidl = 22.4408345339434 pbgidl = -5.46070779382105e-6
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.0678392589988217 lkt1 = -1.08098220053745e-07 wkt1 = -1.1762176426676e-07 pkt1 = 2.86218448731447e-14
+ kt2 = 0.235996541485714 lkt2 = -6.17077285080507e-08 wkt2 = -2.64697796016969e-23
+ at = 392704.922449648 lat = -0.0793644264910523 wat = -0.273858115484662 pat = 6.66400861058066e-8
+ ute = 0.608999778686825 lute = -1.93276019406095e-07 wute = -6.38637550815321e-07 pute = 1.55404784340299e-13
+ ua1 = 1.15501047585414e-09 lua1 = -1.83104660653394e-16 wua1 = -1.14202526933424e-16 pua1 = 2.77898144989255e-23
+ ub1 = -1.27707448617462e-19 lub1 = 1.37901457131676e-25 wub1 = 5.04223532089289e-25 pub1 = -1.22696745851543e-31
+ uc1 = 1.99309798377342e-10 luc1 = -4.83603756466256e-17 wuc1 = -1.77638117517771e-16 puc1 = 4.32261042405393e-23
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.89 pmos
* DC IV MOS Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 6.4e-07 wmax = 8.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.006443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.18282950331546+0*(0.007356/sqrt(l*w*mult))} lvth0 = -1.52767356392756e-07 wvth0 = -4.81927361235598e-07 pvth0 = 8.6627619423399e-14
+ k1 = 2.87836403960321 lk1 = -2.15835788012492e-07 wk1 = -2.4585434495837e-06 pk1 = 3.48345952476648e-13
+ k2 = 0.332552009490551 lk2 = -9.93333847641458e-08 wk2 = -8.51286887496057e-08 pk2 = 1.98944414406093e-14
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -115654.30229193 lvsat = -0.00430554846683723 wvsat = 0.273694675167753 pvsat = -1.62617383445883e-8
+ ua = -1.13210934489676e-08 lua = 1.17505946396009e-15 wua = 1.06916540095196e-14 pua = -1.49484028463845e-21
+ ub = -2.41049583718624e-18 lub = 7.34679397357211e-25 wub = 1.48312809221368e-24 pub = -1.97489777895946e-31
+ uc = 3.47186449884522e-12 luc = -4.70156804581691e-19 wuc = -2.56751950905138e-18 puc = 3.63254106313515e-25
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = -0.0497138271649233 lu0 = 7.33915544591486e-09 wu0 = 5.26251830499949e-08 pu0 = -7.44632089008105e-15
+ a0 = -2.80402064513642 la0 = 5.46713443580799e-07 wa0 = 3.63093322898825e-06 pa0 = -5.15715656781089e-13
+ keta = -2.56245585355066 lketa = 4.28994291474924e-07 wketa = 2.0085560445651e-06 pketa = -3.30472705290292e-13
+ a1 = 0.0
+ a2 = -0.445070893740173 la2 = 2.07061902766929e-07 wa2 = -3.22323651831565e-07 pa2 = 4.62012276062329e-14
+ ags = 15.5143119325553 lags = -2.47254730176527e-06 wags = -9.83869789384694e-06 pags = 1.70542021552364e-12
+ b0 = 1.43374979148345e-05 lb0 = -2.48493431722792e-12 wb0 = -1.27566769372403e-11 pb0 = 2.21095092626587e-18
+ b1 = 1.61347698406525e-07 lb1 = -2.8012782434042e-14 wb1 = -1.43557856145158e-13 pb1 = 2.49241546709859e-20
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-3.81298006685357+0*(0.0/sqrt(l*w*mult))} lvoff = 5.29312077260209e-07 wvoff = 2.83835366085893e-06 pvoff = -4.52578638091009e-13
+ nfactor = {-47.2436340978837+0*(0.1/sqrt(l*w*mult))} lnfactor = 7.30134576688018e-06 wnfactor = 3.90607490409127e-05 pnfactor = -5.38082319552591e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.170367210218553 leta0 = 5.95349459060933e-08 weta0 = -7.72138118459316e-07 peta0 = 8.71937434194953e-14
+ etab = 2.04177785855811 letab = -3.19135830065659e-07 wetab = -1.80239839608268e-06 petab = 2.76610674960542e-13
+ dsub = 0.560954466898676 ldsub = -4.55091431096207e-08 wdsub = -2.18998851535904e-07 pdsub = 3.35003753978878e-14
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.12056326969416 lpclm = -8.87570992562366e-08 wpclm = 9.87921727200869e-07 ppclm = -1.69155827163968e-13
+ pdiblc1 = 0.28884401393627 lpdiblc1 = -3.37875017307465e-08 wpdiblc1 = 4.42765091483021e-07 ppdiblc1 = -6.77533803360373e-14
+ pdiblc2 = -0.013480476217546 lpdiblc2 = 2.10018107759398e-09 wpdiblc2 = 2.2066668515901e-08 ppdiblc2 = -3.25755503382498e-15
+ pdiblcb = -2.02861020764183 lpdiblcb = 2.93803894109094e-07 wpdiblcb = 1.41947856275986e-06 ppdiblcb = -2.06161549605241e-13
+ drout = 1.0
+ pscbe1 = 1457401859.61655 lpscbe1 = -113.952723542214 wpscbe1 = -453.330007749055 ppscbe1 = 7.85793168832055e-5
+ pscbe2 = 1.83190157256176e-07 lpscbe2 = -2.5111972721729e-14 wpscbe2 = -1.52143942285583e-13 ppscbe2 = 2.19107259662728e-20
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 31.8017729021218 lbeta0 = -3.73962829097259e-06 wbeta0 = -1.39614869015835e-05 pbeta0 = 2.19871027693247e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -6.57054687871976e-08 lagidl = 8.70724282637701e-15 wagidl = 5.80339228614216e-14 pagidl = -7.65776249741889e-21
+ bgidl = 1075915243.7619 lbgidl = -10.8815392103429 wbgidl = -52.3619472458668 pbgidl = 7.50545679432816e-6
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.604058755002754 lkt1 = -1.51510050554153e-08 wkt1 = 2.74450783289105e-07 pkt1 = -3.93392263750941e-14
+ kt2 = -0.12
+ at = -136292.704278069 lat = 0.0123309641306765 wat = 0.335579971524386 pat = -3.89986930201676e-8
+ ute = -1.40013053483571 lute = 1.54982610879275e-07 wute = 1.03757183754526e-06 pute = -1.35145998619348e-13
+ ua1 = 1.16054941680031e-09 lua1 = -1.84064769599121e-16 wua1 = -7.16395182317985e-16 pua1 = 1.32172684997975e-22
+ ub1 = 2.09620272744075e-18 lub1 = -2.47586684965903e-25 wub1 = -1.17652157487501e-24 pub1 = 1.68640249499435e-31
+ uc1 = -4.98450921116467e-10 luc1 = 7.25880719489922e-17 wuc1 = 4.144889408748e-16 puc1 = -5.9412015807112e-23
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.90 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 5.5e-07 wmax = 6.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.004443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.0168761+0*(0.005856/sqrt(l*w*mult))}
+ k1 = 0.47866595
+ k2 = -0.0041430645
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 24491.02
+ ua = -9.0913219e-10
+ ub = 1.39839665e-18
+ uc = -6.8009552e-11
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0102961633
+ a0 = 1.2509318
+ keta = 0.0074076058
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.23496304
+ b0 = -2.1309e-8
+ b1 = 2.2477e-9
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.34840646+0*(0.0/sqrt(l*w*mult))}
+ nfactor = {2.0716757+0*(0.1/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.0017402344
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00083787503
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 790097310.0
+ pscbe2 = 9.5178184e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 3.0
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.1731672e-9
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.52561
+ kt2 = -0.052484
+ at = 10000.0
+ ute = -1.2595
+ ua1 = -2.5605e-10
+ ub1 = 4.9434e-19
+ uc1 = 8.1951e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.91 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 5.5e-07 wmax = 6.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.004443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.0168761+0*(0.005856/sqrt(l*w*mult))}
+ k1 = 0.47866595
+ k2 = -0.0041430645
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 24491.02
+ ua = -9.0913219e-10
+ ub = 1.39839665e-18
+ uc = -6.8009552e-11
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0102961633
+ a0 = 1.2509318
+ keta = 0.0074076058
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.23496304
+ b0 = -2.1309e-8
+ b1 = 2.2477e-9
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.34840646+0*(0.0/sqrt(l*w*mult))}
+ nfactor = {2.0716757+0*(0.1/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.0017402344
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00083787503
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 790097310.0
+ pscbe2 = 9.5178184e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 3.0
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.1731672e-9
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.52561
+ kt2 = -0.052484
+ at = 10000.0
+ ute = -1.2595
+ ua1 = -2.5605e-10
+ ub1 = 4.9434e-19
+ uc1 = 8.1951e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.92 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 5.5e-07 wmax = 6.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.004443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.08925744775245+0*(0.005856/sqrt(l*w*mult))} lvth0 = 5.78568577480867e-7
+ k1 = 0.494917388074975 lk1 = -1.29903237519343e-7
+ k2 = -0.0325572332526668 lk2 = 2.27124054829104e-07 pk2 = 5.04870979341448e-29
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 13069.09495219 lvsat = 0.0912993075178117
+ ua = -9.66291472397079e-10 lua = 4.56893464037314e-16
+ ub = 2.21949209410947e-18 lub = -6.56329341502712e-24
+ uc = -6.33446214035016e-11 luc = -3.72883670043541e-17
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0142698174381638 lu0 = -3.17627606214424e-8
+ a0 = 1.2538974524657 la0 = -2.37054625488884e-8
+ keta = 0.00418131295504559 lketa = 2.57888491967021e-8
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.235883554325725 lags = -7.35798213936272e-9
+ b0 = -1.351101479895e-07 lb0 = 9.09651040668094e-13 wb0 = -2.52435489670724e-29
+ b1 = 4.795080260235e-09 lb1 = -2.03620714345863e-14 pb1 = -1.20370621524202e-35
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.444837635940725+0*(0.0/sqrt(l*w*mult))} lvoff = 7.70806983031682e-07 wvoff = -4.2351647362715e-22
+ nfactor = {2.46027311128664+0*(0.1/sqrt(l*w*mult))} lnfactor = -3.10619045433921e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.395686193228354 lpclm = 3.17676376616597e-06 wpclm = 3.30872245021211e-24 ppclm = 3.91275008989622e-28
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00124507074413753 lpdiblc2 = -3.2548529752527e-9
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 780211112.930193 lpscbe1 = 79.0237147135631
+ pscbe2 = 9.45640285822898e-09 lpscbe2 = 4.90915183828849e-16
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.78586633607361e-10 lalpha0 = -6.28169524705797e-16
+ alpha1 = 1.99833416432488e-10 lalpha1 = -7.98002241239631e-16
+ beta0 = -17.6314320251595 lbeta0 = 0.000164914009601124 wbeta0 = -6.7762635780344e-21
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 2.2445470400284e-09 lagidl = -8.56390118773294e-15
+ bgidl = 678903777.929449 lbgidl = 2566.63063353298
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.658049054769999 lkt1 = 1.05863012917712e-6
+ kt2 = -0.046450399725723 lkt2 = -4.82286063491885e-8
+ at = -42713.0729128486 lat = 0.421353408811043 pat = 1.05879118406788e-22
+ ute = -2.153658294925 lute = 7.14730947683921e-6
+ ua1 = -8.85759469220001e-10 lua1 = 5.03348062927607e-15
+ ub1 = 5.65236484917219e-19 lub1 = -5.6669956695524e-25
+ uc1 = 6.07016774048686e-11 luc1 = -4.19702820420277e-16 wuc1 = -1.23259516440783e-32 puc1 = 1.41059322098675e-37
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.93 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 5.5e-07 wmax = 6.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.004443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.871079958408998+0*(0.005856/sqrt(l*w*mult))} lvth0 = -2.92687881458923e-7
+ k1 = 0.475299486095559 lk1 = -5.15623240646724e-8
+ k2 = 0.040644405681078 lk2 = -6.51948315872987e-8
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 39559.583135983 lvsat = -0.0144861655850803
+ ua = -1.08251348411575e-09 lua = 9.21007239869922e-16
+ ub = -8.03800002780308e-20 lub = 2.62087321463009e-24
+ uc = -7.89241966365168e-11 luc = 2.4926142797506e-17
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.00125238287902001 lu0 = 2.02202554661001e-8
+ a0 = 1.3338353970428 la0 = -3.42924694270506e-7
+ keta = 0.0265304661513564 lketa = -6.34588735299472e-8
+ a1 = 0.0
+ a2 = 0.8
+ ags = -0.101537512133451 lags = 1.34007838455259e-6
+ b0 = 2.0447836173e-07 lb0 = -4.46440659558155e-13 pb0 = -1.92592994438724e-34
+ b1 = -9.64701613619999e-10 lb1 = 2.63868439399006e-15 wb1 = -3.94430452610506e-31
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1977606647864+0*(0.0/sqrt(l*w*mult))} lvoff = -2.15854874803786e-7
+ nfactor = {1.14967055274+0*(0.1/sqrt(l*w*mult))} lnfactor = 2.12748854560234e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.1592351855 leta0 = -3.16412877194199e-7
+ etab = -0.1392684955 letab = 2.76612515282979e-7
+ dsub = 0.859000699999999 ldsub = -1.1940108573366e-6
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.498660454442519 lpclm = -3.94664687150745e-07 wpclm = 4.2351647362715e-22
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00057063114206935 lpdiblc2 = -5.61587683608933e-10
+ pdiblcb = -0.424333799999999 lpdiblcb = 7.960072382244e-7
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 9.63030196631712e-09 lpscbe2 = -2.03522732665583e-16
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.87910516027147e-11 lalpha0 = -6.99185148545254e-17 walpha0 = -2.46519032881566e-32 palpha0 = 4.70197740328915e-38
+ alpha1 = 5.73670036880007e-16 lalpha1 = -2.15658830957128e-21 walpha1 = 9.4039548065783e-38 palpha1 = -6.27781712017518e-43
+ beta0 = 44.262864050319 lbeta0 = -8.22508349003348e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -1.5111712326491e-10 lagidl = 1.00279555078445e-15
+ bgidl = 1642192444.1411 lbgidl = -1280.10660221933
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.29548101427894 lkt1 = -3.89226604501367e-7
+ kt2 = -0.0595514414067929 lkt2 = 4.08828123541189e-9
+ at = 85592.4759078148 lat = -0.0910140149053682
+ ute = 0.23572003740572 lute = -2.39428581403369e-6
+ ua1 = 7.57014667690222e-10 lua1 = -1.52667175706473e-15
+ ub1 = 3.3072320827312e-19 lub1 = 3.69791212172155e-25
+ uc1 = -1.34630329173249e-10 luc1 = 3.6032390406437e-16 wuc1 = 4.93038065763132e-32
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.94 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 5.5e-07 wmax = 6.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.004443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.049504128414+0*(0.005856/sqrt(l*w*mult))} lvth0 = 6.29717967305065e-8
+ k1 = 0.414136178847399 lk1 = 7.03568204787615e-8
+ k2 = 0.019004695517398 lk2 = -2.20595750090491e-08 wk2 = -1.32348898008484e-23
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -120709.932052356 lvsat = 0.304985149281413 pvsat = 5.29395592033938e-23
+ ua = -2.38835009088599e-10 lua = -7.60729124183748e-16
+ ub = 1.22011089563328e-18 lub = 2.85552931560295e-26
+ uc = -1.0751845924825e-10 luc = 8.1924173043452e-17
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0140859613026 lu0 = -5.3614040816021e-09 wu0 = -1.32348898008484e-23
+ a0 = 1.1025970552 la0 = 1.18011479581738e-7
+ keta = -0.0111645336712126 lketa = 1.16800020263728e-8
+ a1 = 0.0
+ a2 = 1.1973352 la2 = -7.920233528976e-7
+ ags = 0.68894229203862 lags = -2.35615047336159e-7
+ b0 = -1.61612814364e-07 lb0 = 2.83302793214707e-13 pb0 = -7.22223729145213e-35
+ b1 = 2.8206905647e-09 lb1 = -4.90688167995797e-15 wb1 = 7.88860905221012e-31 pb1 = 3.76158192263132e-37
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.35231008046714+0*(0.0/sqrt(l*w*mult))} lvoff = 9.22143483504274e-8
+ nfactor = {-0.341843953883803+0*(0.1/sqrt(l*w*mult))} lnfactor = 5.10058108920683e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = -0.485738951 leta0 = 9.69238578108438e-07 weta0 = -1.57164316385075e-22 peta0 = -2.20881053461883e-29
+ etab = 0.162904101 letab = -3.25719603879139e-07 wetab = 5.12851979782877e-23 petab = 2.20881053461883e-29
+ dsub = 0.26
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.0742494148848616 lpclm = 7.47338325954558e-7
+ pdiblc1 = 0.389494937293899 lpdiblc1 = 1.00676068445305e-9
+ pdiblc2 = 0.000148737715861299 lpdiblc2 = 2.79388514801769e-10
+ pdiblcb = 0.1736676 lpdiblcb = -3.960116764488e-07 ppdiblcb = -1.51461293802434e-28
+ drout = 0.233817461872679 ldrout = 6.50192048185637e-7
+ pscbe1 = 801195690.883978 lpscbe1 = -2.38341607528855
+ pscbe2 = 1.00453763670072e-08 lpscbe2 = -1.03090630838839e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -9.19286376348734e-11 lalpha0 = 1.9065000905095e-16 walpha0 = -6.16297582203915e-33 palpha0 = -5.87747175411144e-39
+ alpha1 = -9.93348130700257e-11 lalpha1 = 1.98006844545353e-16 walpha1 = -5.91922531345265e-33 palpha1 = 8.26497941477509e-38
+ beta0 = -1.89174393923941 lbeta0 = 9.75089908035558e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 7.57762120486598e-11 lagidl = 5.50520443557167e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.46303225874108 lkt1 = -5.52403419676924e-8
+ kt2 = -0.0552956877620159 lkt2 = -4.39487422336052e-9
+ at = 7282.96884286986 lat = 0.0650833012884552
+ ute = -1.74526153944298 lute = 1.55448004039875e-6
+ ua1 = -1.01421246704804e-09 lua1 = 2.00398259724017e-15 wua1 = -7.39557098644699e-32 pua1 = -3.76158192263132e-37
+ ub1 = 1.51236168895956e-18 lub1 = -1.98561367364239e-24 wub1 = -7.3468396926393e-40
+ uc1 = 9.45390689071462e-11 luc1 = -9.64881655664091e-17 puc1 = 4.70197740328915e-38
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.95 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 5.5e-07 wmax = 6.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.004443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.021185345124+0*(0.005856/sqrt(l*w*mult))} lvth0 = 3.48416731747835e-8
+ k1 = 0.433942827763722 lk1 = 5.06821234575217e-8
+ k2 = 0.0053098971143308 lk2 = -8.45601135294313e-09 pk2 = -3.15544362088405e-30
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 281821.671312781 lvsat = -0.0948647885421043
+ ua = -2.19856609529999e-10 lua = -7.79581089644489e-16
+ ub = 6.40974805810801e-19 lub = 6.03833178348113e-25
+ uc = -3.68425960659401e-11 luc = 1.17191524616627e-17
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0119524255404 lu0 = -3.24208193464985e-9
+ a0 = 1.3370384272 la0 = -1.14868043997993e-7
+ keta = 0.0102543614029353 lketa = -9.59620036879108e-09 wketa = 1.65436122510606e-24 pketa = -1.57772181044202e-30
+ a1 = 0.0
+ a2 = 0.00532960000000049 la2 = 3.920411057952e-7
+ ags = 0.0750739951768802 lags = 3.74163658931889e-7
+ b0 = 2.21467272524e-07 lb0 = -9.72252141344452e-14
+ b1 = -2.05039325756e-08 lb1 = 1.82623528209814e-14 wb1 = 3.15544362088405e-30 pb1 = 3.00926553810506e-36
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.17299845369812+0*(0.0/sqrt(l*w*mult))} lvoff = -8.59027043610566e-8
+ nfactor = {7.20701764227201+0*(0.1/sqrt(l*w*mult))} lnfactor = -2.39798999099538e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.49
+ etab = -0.327795373275 letab = 1.61710830498242e-7
+ dsub = 0.22285388835452 ldsub = 3.68986442496979e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.724860464581081 lpclm = -4.64478834943812e-8
+ pdiblc1 = 0.582254436329561 lpdiblc1 = -1.90468574568633e-07 wpdiblc1 = 4.2351647362715e-22
+ pdiblc2 = -6.97233132010396e-05 lpdiblc2 = 4.96394156488494e-10
+ pdiblcb = -0.225
+ drout = 0.940647677979241 ldrout = -5.19292650212225e-8
+ pscbe1 = 797608618.23204 lpscbe1 = 1.17975949864194
+ pscbe2 = 1.69084195225236e-08 lpscbe2 = -7.84822787040275e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 6.80525548816681 lbeta0 = 1.11183906313476e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 9.2751125890816e-10 lagidl = -2.95540344420154e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.527763005202081 lkt1 = 9.05916826038275e-9
+ kt2 = -0.0440516586270121 lkt2 = -1.55639956362672e-8
+ at = 79613.5535857882 lat = -0.00676541709890555
+ ute = -0.267515207816925 lute = 8.65784548339858e-8
+ ua1 = 1.6847864446152e-09 lua1 = -6.77035583673575e-16
+ ub1 = -1.43727939498936e-18 lub1 = 9.44376901405261e-25 pub1 = -3.50324616081204e-46
+ uc1 = -2.91537921926444e-11 luc1 = 2.63806536927348e-17 wuc1 = 6.16297582203915e-33 puc1 = 1.0285575569695e-38
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.96 pmos
* DC IV MOS Parameters
+ lmin = 2.5e-07 lmax = 5e-07 wmin = 5.5e-07 wmax = 6.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.006443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.939594243016002+0*(0.007356/sqrt(l*w*mult))} lvth0 = -5.41031795697235e-9
+ k1 = 0.494267157497442 lk1 = 2.09218392753482e-8
+ k2 = -0.00919181642799757 lk2 = -1.30176499739792e-9
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 67329.9919879199 lvsat = 0.0109521075526635
+ ua = -2.0449807407592e-09 lua = 1.20821999007862e-16
+ ub = 2.041231234016e-18 lub = -8.69665274297851e-26
+ uc = -2.58807559379872e-11 luc = 6.31126017661872e-18
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.00522382485816002 lu0 = 7.73924687250611e-11
+ a0 = 1.38850638568 la0 = -1.402591436986e-7
+ keta = -0.008445362407908 lketa = -3.7091602339729e-10
+ a1 = 0.0
+ a2 = 1.06891451743248 la2 = -1.32665750201105e-7
+ ags = 1.23423871552472 lags = -1.97696345875074e-7
+ b0 = 4.8132028632e-08 lb0 = -1.17123515832536e-14
+ b1 = 3.2587934928e-08 lb1 = -7.92988290950966e-15
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.2740601181368+0*(0.0/sqrt(l*w*mult))} lvoff = -3.60451449502073e-8
+ nfactor = {1.68816362963119+0*(0.1/sqrt(l*w*mult))} lnfactor = 3.24670409892803e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.49
+ etab = 4.850105e-05 letab = -2.70107735049e-11 petab = 3.08148791101958e-33
+ dsub = -0.023901594981119 ldsub = 1.58632500887536e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.624438894129922 lpclm = 3.09389322885369e-9
+ pdiblc1 = -0.0625215999738398 lpdiblc1 = 1.27623945629214e-07 ppdiblc1 = -5.04870979341448e-29
+ pdiblc2 = -0.0089245210323659 lpdiblc2 = 4.86480235366586e-09 wpdiblc2 = 1.65436122510606e-24 ppdiblc2 = -7.88860905221012e-31
+ pdiblcb = -0.225
+ drout = 1.22833572426512 ldrout = -1.93856710399806e-07 wdrout = 8.470329472543e-22
+ pscbe1 = 800069244.26128 lpscbe1 = -0.0341608253716004
+ pscbe2 = -6.99090056320879e-09 lpscbe2 = 3.9422149020523e-15 ppscbe2 = -1.1284745767894e-36
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.83100208558321 lbeta0 = 1.12461288258562e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 5.5080962010832e-10 lagidl = -1.09699111337918e-16
+ bgidl = 730034204.006401 lbgidl = 133.18438586389
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.50680115016 lkt1 = -1.28211138236603e-9
+ kt2 = -0.132062202816 lkt2 = 2.78549502128398e-8
+ at = 65261.4810880001 lat = 0.000315005643008265
+ ute = -0.0012549260000001 lute = -4.47778600770119e-8
+ ua1 = 2.2472125128e-10 lua1 = 4.32700586760273e-17
+ ub1 = 5.1394790896e-19 lub1 = -1.82376742705086e-26
+ uc1 = 4.74348323563201e-11 luc1 = -1.14034251650022e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.24e-6
+ sbref = 1.24e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.97 pmos
* DC IV MOS Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 5.5e-07 wmax = 6.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.006443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.772463663771422+0*(0.007356/sqrt(l*w*mult))} lvth0 = -4.60795388491882e-8
+ k1 = -0.41547953916943 lk1 = 2.4229778094887e-7
+ k2 = 0.438589349394086 lk2 = -1.10263938326212e-07 wk2 = 5.29395592033938e-23 pk2 = 4.41762106923767e-29
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 92623.7868717136 lvsat = 0.00479716609323066
+ ua = -1.55915274021428e-09 lua = 2.60158501126276e-18
+ ub = 9.27892317999923e-20 lub = 3.87163452505452e-25
+ uc = 6.09622494694269e-15 luc = 1.20053449946549e-20
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.00281915098371424 lu0 = 6.62540999984932e-10
+ a0 = -0.397764477428577 la0 = 2.94408435588514e-7
+ keta = -0.184161871607297 lketa = 4.23875878921637e-08 wketa = 2.64697796016969e-23 pketa = -6.31088724176809e-30
+ a1 = 0.0
+ a2 = 0.164955374457998 la2 = 8.73018597320191e-8
+ ags = -1.62902379023886 lags = 4.99044225752424e-07 pags = 2.01948391736579e-28
+ b0 = 1.23812857142857e-09 lb0 = -3.01283730314285e-16
+ b1 = -1.86798933828571e-10 lb1 = 4.54552789599769e-17
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.403685441391142+0*(0.0/sqrt(l*w*mult))} lvoff = -4.50237804014223e-9
+ nfactor = {-5.5978371627743+0*(0.1/sqrt(l*w*mult))} lnfactor = 2.09763127071517e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 1.39713389074943 leta0 = -2.20740146707184e-7
+ etab = 0.244655617911143 letab = -5.95492173762616e-08 wetab = 1.6130021944784e-23 petab = -1.1339875512552e-29
+ dsub = 1.53653693089571 ldsub = -2.21081489122281e-07 pdsub = 2.01948391736579e-28
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.664807054980852 lpclm = -6.72921429629145e-9
+ pdiblc1 = 1.18699067550629 lpdiblc1 = -1.76429872461569e-7
+ pdiblc2 = 0.0300992129326342 lpdiblc2 = -4.63115502190936e-09 wpdiblc2 = -2.64697796016969e-23
+ pdiblcb = -0.78214353300956 lpdiblcb = 1.35574193035481e-7
+ drout = -0.975627884694001 ldrout = 3.42451386277088e-7
+ pscbe1 = 799752699.066856 lpscbe1 = 0.0428666491488912
+ pscbe2 = 2.95389305828886e-08 lpscbe2 = -4.94688114937674e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 11.56376242988 lbeta0 = -5.52523148401942e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -1.10815918728486e-08 lagidl = 2.72090620315522e-15 wagidl = 2.76101316827354e-30 pagidl = 4.70197740328915e-37
+ bgidl = 1964163557.12 lbgidl = -167.126182664067
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.238369297999997 lkt1 = -6.66017814232763e-8
+ kt2 = 0.235996541485714 lkt2 = -6.17077285080508e-08 wkt2 = -5.29395592033938e-23 pkt2 = -2.52435489670724e-29
+ at = -4339.24200000009 lat = 0.017251506397796
+ ute = -0.316907829714285 lute = 3.20324862070149e-8
+ ua1 = 9.8943770542857e-10 lua1 = -1.42814513843578e-16 wua1 = 7.88860905221012e-31
+ ub1 = 6.03324423999999e-19 lub1 = -3.9986376687312e-26
+ uc1 = -5.82329727011429e-11 luc1 = 1.43095671820707e-17 wuc1 = -2.31111593326468e-32 puc1 = 3.67341984631965e-40
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.98 pmos
* DC IV MOS Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 5.5e-07 wmax = 6.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.006443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.520352091175162+0*(0.007356/sqrt(l*w*mult))} lvth0 = -8.97800546198801e-08 wvth0 = -2.49123788935557e-07 pvth0 = 4.31826193265113e-14
+ k1 = -4.11333191723232 lk1 = 8.83276116457536e-07 wk1 = 2.36392430141515e-06 pk1 = -4.097579105587e-13
+ k2 = 1.33266162872819 lk2 = -2.65240639081427e-07 wk2 = -7.74946497763736e-07 pk2 = 1.3432767602937e-13
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 553155.212815385 lvsat = -0.0750304302169931 wvsat = -0.187611471163299 pvsat = 3.25201971885039e-8
+ ua = 1.02679182791027e-08 lua = -2.04747925133511e-15 wua = -4.19919843562542e-15 pua = 7.27880658434437e-22
+ ub = -4.24535660405064e-18 lub = 1.13912897540013e-24 wub = 2.74870899424445e-24 pub = -4.76455719644343e-31
+ uc = 2.07223916932761e-13 luc = -2.2857726878783e-20 wuc = -3.15759131873796e-19 puc = 5.47330564007401e-26
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0444091931970076 lu0 = -6.5465937371829e-09 wu0 = -1.22954360850881e-08 pu0 = 2.13126630011701e-15
+ a0 = -10.6730705149987 la0 = 2.07550943352884e-06 wa0 = 9.05854899813677e-06 pa0 = -1.57019076623903e-12
+ keta = -0.441264945469912 lketa = 8.69533205093617e-08 wketa = 5.45481161005485e-07 pketa = -9.45526134863688e-14
+ a1 = 0.0
+ a2 = -7.2643021704831 la2 = 1.37507450405702e-06 wa2 = 4.38118793129792e-06 pa2 = -7.59426353635319e-13
+ ags = 21.1495017276852 lags = -3.4493398304735e-06 wags = -1.37255261005574e-05 pags = 2.37915524321842e-12
+ b0 = -1.01826005104488e-05 lb0 = 1.76494493828017e-12 wb0 = 4.15586969483117e-12 pb0 = -7.20370141162646e-19
+ b1 = 3.81162611686897e-07 lb1 = -6.60568888592154e-14 wb1 = -2.95173478023971e-13 pb1 = 5.11647803337191e-20
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {4.55595098084441+0*(0.0/sqrt(l*w*mult))} lvoff = -8.64195836197608e-07 wvoff = -2.93405125162859e-06 pvoff = 5.08582575854796e-13
+ nfactor = {8.69002721260188+0*(0.1/sqrt(l*w*mult))} lnfactor = -3.78998564383784e-07 wnfactor = 4.80942434563544e-07 pnfactor = -8.33655997223732e-14
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = -6.31559897469831 leta0 = 1.1161695427238e-06 weta0 = 3.70150646705085e-06 peta0 = -6.4161172798566e-13
+ etab = -1.28158713182753 letab = 2.05006648377941e-07 wetab = 4.89866683788896e-07 petab = -8.49125112345996e-14
+ dsub = 0.0907377406737719 ldsub = 2.95304509124099e-08 wdsub = 1.0532946768726e-07 pdsub = -1.82575992699743e-14
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 15.1235848598275 lpclm = -2.5129848414328e-06 wpclm = -8.6705531910252e-06 ppclm = 1.50293634902593e-12
+ pdiblc1 = 6.28425096755649 lpdiblc1 = -1.05997877696497e-06 wpdiblc1 = -3.69252009060229e-06 ppdiblc1 = 6.4005404746482e-13
+ pdiblc2 = 0.127385736727115 lpdiblc2 = -2.1494606483397e-08 wpdiblc2 = -7.5094703106218e-08 ppdiblc2 = 1.30167656470256e-14
+ pdiblcb = -2.16260086989224 lpdiblcb = 3.7485990689605e-07 wpdiblcb = 1.51189757691991e-06 ppdiblcb = -2.62069302188144e-13
+ drout = 1.0
+ pscbe1 = 801197746.521767 lpscbe1 = -0.207614986587942 wpscbe1 = -0.718339133996778 ppscbe1 = 1.24515468808914e-7
+ pscbe2 = -2.57115376447668e-08 lpscbe2 = 4.6301245122686e-15 wpscbe2 = -8.0556276608785e-15 ppscbe2 = 1.39634638748135e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 13.1646409435277 lbeta0 = -8.30016228200577e-07 wbeta0 = -1.10667050277243e-06 pbeta0 = 1.91828051609566e-13
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.17461625048231e-08 lagidl = -1.23601108516162e-15 wagidl = 4.61226430047438e-15 pagidl = -7.99480669315629e-22
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = 1.93948854361926 lkt1 = -4.44107303973876e-07 wkt1 = -1.4799411262665e-06 pkt1 = 2.56530034944782e-13
+ kt2 = -0.12
+ at = 886727.42584506 lat = -0.137204207673131 wat = -0.370040183671028 pat = 6.41420253571686e-8
+ ute = 5.88488445721897 lute = -1.04297378522542e-06 wute = -3.98721043010752e-06 pute = 6.91135081533978e-13
+ ua1 = -6.25358620211367e-10 lua1 = 1.37091051650198e-16 wua1 = 5.15420956128132e-16 pua1 = -8.9342037693338e-23
+ ub1 = 5.09221917644162e-19 lub1 = -2.36748364406034e-26 wub1 = -8.19139397681272e-26 pub1 = 1.41987984915277e-32
+ uc1 = 6.3301884706147e-10 luc1 = -1.05510640751941e-16 wuc1 = -3.65933506261741e-16 puc1 = 6.34301821083976e-23
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.99 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 4.2e-07 wmax = 5.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.004443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.13181153747554+0*(0.005856/sqrt(l*w*mult))} wvth0 = 6.89316321295417e-8
+ k1 = 0.5536725055272 wk1 = -4.49845966263051e-8
+ k2 = -0.0764006435052808 wk2 = 4.33359193993009e-8
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -248939.518899277 wvsat = 0.163987832946638
+ ua = -1.34314287141275e-09 wua = 2.60294520893984e-16
+ ub = 4.39741842647386e-18 wub = -1.79863991807034e-24
+ uc = -4.87091391354924e-12 wuc = -3.78669057109717e-17
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.022432676439988 wu0 = -7.27877909090531e-9
+ a0 = 0.0081446176441542 wa0 = 7.45351918877897e-7
+ keta = -0.0550604796320326 wketa = 3.74647469867952e-8
+ a1 = 0.0
+ a2 = 0.0791263930769226 wa2 = 4.32338322937981e-7
+ ags = 0.592480648626646 wags = -2.14418397136484e-7
+ b0 = -6.29827212832308e-08 wb0 = 2.49934892845916e-14
+ b1 = 1.41734032646154e-09 wb1 = 4.98001737399239e-16
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.425953345210784+0*(0.0/sqrt(l*w*mult))} wvoff = 4.65081395394634e-8
+ nfactor = {3.15617132384077+0*(0.1/sqrt(l*w*mult))} wnfactor = -6.50417791332635e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.00752026452741314 wpclm = -3.46652798468104e-9
+ pdiblc1 = 0.39
+ pdiblc2 = -0.00486236335036257 wpdiblc2 = 3.41867350676308e-9
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 1313834677.59128 wpscbe1 = -314.107401061401
+ pscbe2 = 8.13931185585953e-09 wpscbe2 = 8.26748547497198e-16
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 4.61340153846154e-10 walpha0 = -2.16710938816031e-16
+ alpha1 = 4.61340153846154e-10 walpha1 = -2.16710938816031e-16
+ beta0 = -94.5618415384615 wbeta0 = 5.85119534803283e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 3.37464993751129e-09 wagidl = -1.32032210025704e-15
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -1.20164129383077 wkt1 = 4.05444495430912e-7
+ kt2 = -0.0291177113072416 wkt2 = -1.40137493864301e-8
+ at = -261141.0696175 wat = 0.162614741602753
+ ute = -4.72388485901538 wute = 2.07773779699258e-6
+ ua1 = -3.41965361665512e-09 wua1 = 1.8973465929807e-15
+ ub1 = 1.39510181602126e-18 wub1 = -5.40224873216586e-25
+ uc1 = -2.12165063617345e-10 wuc1 = 1.32159289320226e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.100 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 4.2e-07 wmax = 5.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.004443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.097385963809+0*(0.005856/sqrt(l*w*mult))} lvth0 = -6.8828213015911e-07 wvth0 = 4.82851628425066e-08 pvth0 = 4.12791838962311e-13
+ k1 = 0.578425765536448 lk1 = -4.94900293966763e-07 wk1 = -5.98301712414229e-08 pk1 = 2.96812591084273e-13
+ k2 = -0.062650490227771 lk2 = -2.7491146202906e-07 wk2 = 3.508937222231e-08 pk2 = 1.64876005042525e-13
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -390400.785728908 lvsat = 2.82828292163301 wvsat = 0.248828124329828 pvsat = -1.69624062164261e-6
+ ua = -1.34647393985968e-09 lua = 6.6599177360481e-17 wua = 2.62292303212693e-16 pua = -3.9942337148363e-23
+ ub = 4.36537977955187e-18 lub = 6.40559496973946e-25 wub = -1.77942498948033e-24 pub = -3.84170561946047e-31
+ uc = 6.18083202565629e-12 luc = -2.20961292052666e-16 wuc = -4.4495104134392e-17 puc = 1.32519811410508e-22
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0225016375839453 lu0 = -1.37876346000426e-09 wu0 = -7.32013799909675e-09 pu0 = 8.26902630782492e-16
+ a0 = -0.780226219859202 la0 = 1.57621646235477e-05 wa0 = 1.218171179378e-06 pa0 = -9.45323528808866e-12
+ keta = -0.0903377472911431 lketa = 7.05310336025064e-07 wketa = 5.8622013102659e-08 pketa = -4.23004372610411e-13
+ a1 = 0.0
+ a2 = -0.401055806541017 la2 = 9.60044501854497e-06 wa2 = 7.20323851737685e-07 pa2 = -5.7577920164012e-12
+ ags = 0.80716748652396 lags = -4.29230651423221e-06 wags = -3.43175153608062e-07 pags = 2.57427735191996e-12
+ b0 = 3.03751078259463e-07 lb0 = -7.33223281028131e-12 wb0 = -1.94952246467502e-13 pb0 = 4.3974494365503e-18
+ b1 = -1.17892346664391e-08 lb1 = 2.6404351765541e-13 wb1 = 8.41854207810647e-15 pb1 = -1.58358040174395e-19
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.284051562360231+0*(0.0/sqrt(l*w*mult))} lvoff = -2.83709030733373e-06 wvoff = -3.85963478912499e-08 pvoff = 1.70152278251901e-12
+ nfactor = {3.40491942273428+0*(0.1/sqrt(l*w*mult))} lnfactor = -4.97330481803539e-06 wnfactor = -7.99602523408848e-07 pnfactor = 2.98270077283915e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -2.03464159443462e-06 lcit = 2.4061265710639e-10 wcit = 7.21768242605774e-12 pcit = -1.44305564320832e-16
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.48248108775496 lpclm = -2.94893902755465e-05 wpclm = -8.88062777020979e-07 ppclm = 1.76860318005149e-11
+ pdiblc1 = 0.39
+ pdiblc2 = -0.00947587760059476 lpdiblc2 = 9.22395497727087e-08 wpdiblc2 = 6.18559269292869e-09 ppdiblc2 = -5.53199505076938e-14
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 1656546466.01729 lpscbe1 = -6851.95262258565 wpscbe1 = -519.646123017949 ppscbe1 = 0.00410940514016528
+ pscbe2 = 7.14432644037761e-09 lpscbe2 = 1.98930797168004e-14 wpscbe2 = 1.42348328954624e-15 ppscbe2 = -1.19307193941293e-20
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 7.02032985734846e-10 lalpha0 = -4.8122531421278e-15 walpha0 = -3.61064587337185e-16 palpha0 = 2.88611128641664e-21
+ alpha1 = 7.02032985734846e-10 lalpha1 = -4.8122531421278e-15 walpha1 = -3.61064587337185e-16 palpha1 = 2.88611128641664e-21
+ beta0 = -155.154652694166 lbeta0 = 0.00121145255380617 wbeta0 = 9.4852019347035e-05 pbeta0 = -7.26559219815329e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 4.04976259448444e-09 lagidl = -1.34977555389422e-14 wagidl = -1.72521565039797e-15 pagidl = 8.0951736019874e-21
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -1.32198770977512 lkt1 = 2.4061265710639e-06 wkt1 = 4.77621319691489e-07 pkt1 = -1.44305564320832e-12
+ kt2 = -0.0291177113072416 wkt2 = -1.40137493864301e-8
+ at = -261141.0696175 wat = 0.162614741602753
+ ute = -4.72388485901539 wute = 2.07773779699258e-6
+ ua1 = -3.41965361665512e-09 wua1 = 1.8973465929807e-15
+ ub1 = 1.39510181602126e-18 wub1 = -5.40224873216587e-25
+ uc1 = -2.28532176185776e-10 luc1 = 3.2723321366469e-16 wuc1 = 1.41975337419665e-16 puc1 = -1.96255567476332e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.101 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 4.2e-07 wmax = 5.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.004443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.75153208386546+0*(0.005856/sqrt(l*w*mult))} lvth0 = 4.5405289088408e-06 wvth0 = 3.97194047266617e-07 pvth0 = -2.37615480544253e-12
+ k1 = 0.591486079244702 lk1 = -5.99295795822876e-07 wk1 = -5.79163192932525e-08 pk1 = 2.81514525580591e-13
+ k2 = -0.306675478305555 lk2 = 1.67566274812264e-06 wk2 = 1.64400279348158e-07 pk2 = -8.68749782700989e-13
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -89264.695165759 lvsat = 0.421200365763145 wvsat = 0.061373892419677 pvsat = -1.97855586454384e-7
+ ua = -1.56280940607658e-09 lua = 1.79584168021972e-15 wua = 3.57756977884394e-16 pua = -8.03023748859311e-22
+ ub = 1.05062939588489e-17 lub = -4.84458431671395e-23 wub = -4.9699447813229e-24 pub = 2.51187325299413e-29
+ uc = 5.88486504932358e-14 luc = -1.72026209704606e-16 wuc = -3.80257366178169e-17 puc = 8.08079702043027e-23
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.052594110308384 lu0 = -2.41918069202224e-07 wu0 = -2.29846957194301e-08 pu0 = 1.26039007109917e-13
+ a0 = 1.20536821402319 la0 = -1.09362817392919e-07 wa0 = 2.91050322278374e-08 pa0 = 5.13723304403464e-14
+ keta = -0.0169846600745327 lketa = 1.18974316559218e-07 wketa = 1.26941272299e-08 pketa = -5.58872572040236e-14
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.274428699785491 lags = -3.3945326121706e-08 wags = -2.31171503373601e-08 pags = 1.59455521721278e-14
+ b0 = -1.836440293434e-06 lb0 = 9.77504020834815e-12 wb0 = 1.0203594843552e-12 pb0 = -5.31694800328061e-18
+ b1 = 4.80223568679698e-08 lb1 = -2.14050749797058e-13 wb1 = -2.59252219727314e-14 pb1 = 1.16163274076201e-19
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.35203925379799+0*(0.0/sqrt(l*w*mult))} lvoff = 5.69969629016802e-06 wvoff = 5.44087094137278e-07 pvoff = -2.95606291661842e-12
+ nfactor = {6.14613801227154+0*(0.1/sqrt(l*w*mult))} lnfactor = -2.688479153609e-05 wnfactor = -2.21056872461946e-06 pnfactor = 1.42610305256916e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 2.80670076923077e-05 wcit = -1.08355469408015e-11
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -4.04025260894415 lpclm = 1.46556868461589e-05 wpclm = 2.18580028020751e-06 ppclm = -6.88439458162576e-12
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00394223301804862 lpdiblc2 = -1.50159437234969e-08 wpdiblc2 = -1.61760203591244e-09 ppdiblc2 = 7.05362243975163e-15
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 753729551.529228 lpscbe1 = 364.56812703449 wpscbe1 = 15.8821098940512 ppscbe1 = -0.00017125303404306
+ pscbe2 = 9.34969932120297e-09 lpscbe2 = 2.26478886432963e-15 wpscbe2 = 6.39946140437645e-17 ppscbe2 = -1.06386690366568e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 4.62551696386713e-10 lalpha0 = -2.89799825169237e-15 walpha0 = -1.70305831474426e-16 palpha0 = 1.36131207434613e-21
+ alpha1 = 5.60571636959512e-10 lalpha1 = -3.68150476743067e-15 walpha1 = -2.16349934002962e-16 palpha1 = 1.72935814876337e-21
+ beta0 = -98.7779539734964 lbeta0 = 0.000760814545607688 wbeta0 = 4.86669935956439e-05 pbeta0 = -3.57386698445756e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 7.30384235137417e-09 lagidl = -3.95087149147197e-14 wagidl = -3.0342729004762e-15 pagidl = 1.85589106632132e-20
+ bgidl = -481345804.894464 lbgidl = 11840.8977134035 wbgidl = 695.850637351896 pbgidl = -0.00556216934186913
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -1.69426959642841 lkt1 = 5.38190152236133e-06 wkt1 = 6.21465187339403e-07 pkt1 = -2.59284829654537e-12
+ kt2 = 0.011922586986256 lkt2 = -3.28048975880749e-07 wkt2 = -3.50087434712131e-08 pkt2 = 1.67820084027671e-13
+ at = -580986.793542041 lat = 2.55663497918354 wat = 0.322825465412337 pat = -1.28061846663466e-6
+ ute = -10.1128068191824 lute = 4.30754746832378e-05 wute = 4.77343724606491e-06 pute = -2.1547636842849e-11
+ ua1 = -8.66252479772217e-09 lua1 = 4.19080414407281e-14 wua1 = 4.66405434699961e-15 pua1 = -2.2115230225094e-20
+ ub1 = 3.43513366812909e-18 lub1 = -1.63066641246639e-23 wub1 = -1.72119845043329e-24 pub1 = 9.43992097176223e-30
+ uc1 = -1.23024314965974e-11 luc1 = -1.40116422128962e-15 wuc1 = 4.37836448816047e-17 puc1 = 5.8862381977246e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.102 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 4.2e-07 wmax = 5.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.004443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.244253887818843+0*(0.005856/sqrt(l*w*mult))} lvth0 = -1.47854238800361e-06 wvth0 = -3.75934046593098e-07 pvth0 = 7.1120699063503e-13
+ k1 = 0.420797466108852 lk1 = 8.23215291798104e-08 wk1 = 3.26871613712719e-08 pk1 = -8.02957966893227e-14
+ k2 = 0.221708244813498 lk2 = -4.34352051990156e-07 wk2 = -1.08591625221724e-07 pk2 = 2.21399163510295e-13
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 61722.9094512185 lvsat = -0.181744173282808 wvsat = -0.0132922820836173 pvsat = 1.00311685504252e-7
+ ua = -2.01297051172557e-09 lua = 3.59348712952987e-15 wua = 5.58034344744174e-16 pua = -1.60279896848041e-21
+ ub = -4.21144103905679e-18 lub = 1.03270472739271e-23 wub = 2.47757163573146e-24 pub = -4.62171778390572e-30
+ uc = -5.38300131134682e-11 luc = 4.31702297541683e-17 wuc = -1.5050040833317e-17 puc = -1.09417488483803e-23
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = -0.0273162283959642 lu0 = 7.71909229387209e-08 wu0 = 1.71338017770039e-08 pu0 = -3.41677134454981e-14
+ a0 = 1.54668355629703 la0 = -1.47235034367806e-06 wa0 = -1.27654023297083e-07 pa0 = 6.77364223712119e-13
+ keta = 0.0581517503400803 lketa = -1.81070766333052e-07 wketa = -1.89646185461705e-08 pketa = 7.05368153358982e-14
+ a1 = 0.0
+ a2 = 0.8
+ ags = -0.769227313045396 lags = 4.13372588884437e-06 wags = 4.00441750116493e-07 pags = -1.67546830024846e-12
+ b0 = 1.22393762790181e-06 lb0 = -2.44608323928315e-12 wb0 = -6.11412743104268e-13 pb0 = 1.19927003997794e-18
+ b1 = 1.16548799309345e-08 lb1 = -6.88231221802718e-14 wb1 = -7.56849559861051e-15 pb1 = 4.28586610908223e-20
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {0.315997186170879+0*(0.0/sqrt(l*w*mult))} lvoff = -9.61337010944397e-07 wvoff = -3.0812226380039e-07 pvoff = 4.4709709638967e-13
+ nfactor = {-3.10848396148035+0*(0.1/sqrt(l*w*mult))} lnfactor = 1.00720420673285e-05 wnfactor = 2.55379495629844e-06 pnfactor = -4.76468400713777e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 2.80670076923077e-05 wcit = -1.08355469408015e-11
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.1592351855 leta0 = -3.16412877194199e-7
+ etab = -0.1392684955 letab = 2.76612515282979e-7
+ dsub = 0.8590007 ldsub = -1.1940108573366e-6
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.0251475491022051 lpclm = -1.57883009017358e-06 wpclm = 2.83985671577193e-07 ppclm = 7.10193963972804e-13
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00362348161614442 lpdiblc2 = -1.37430616377196e-08 wpdiblc2 = -1.83092325959283e-09 ppdiblc2 = 7.90548618848105e-15
+ pdiblcb = -1.14460685958738 lpdiblcb = 3.67230101745096e-06 wpdiblcb = 4.31978149357668e-07 ppdiblcb = -1.72503475899965e-12
+ drout = 0.56
+ pscbe1 = 889897293.439555 lpscbe1 = -179.195691110215 wpscbe1 = -53.9152005414844 ppscbe1 = 0.000107471218016962
+ pscbe2 = 1.00279120245314e-08 lpscbe2 = -4.43543695954518e-16 wpscbe2 = -2.3846353105557e-16 ppscbe2 = 1.43950700569001e-22
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -5.4251798649734e-10 lalpha0 = 1.11558470561647e-15 walpha0 = 3.48635561390011e-16 palpha0 = -7.10996309552359e-22
+ alpha1 = -7.21474037069614e-10 lalpha1 = 1.43813694040546e-15 walpha1 = 4.32698770289142e-16 palpha1 = -8.62512705937055e-22
+ beta0 = 277.427250265833 lbeta0 = -0.00074149999227899 wbeta0 = -0.000139838521950542 pbeta0 = 3.95379539994421e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -4.23641794250093e-09 lagidl = 6.57544504670294e-15 wagidl = 2.45012730099042e-15 pagidl = -3.34215306851105e-21
+ bgidl = 3962691609.78892 lbgidl = -5905.64576807343 wbgidl = -1391.70127470379 pbgidl = 0.0027741310355155
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.07695428438333 lkt1 = -1.07658517121012e-06 wkt1 = -1.31059701746399e-07 pkt1 = 4.12237938986756e-13
+ kt2 = -0.0749495632854872 lkt2 = 1.8860882941113e-08 wkt2 = 9.23490349139609e-09 pkt2 = -8.85975264670087e-15
+ at = 201781.238246617 lat = -0.569222347343314 wat = -0.0696833039403501 pat = 2.86801717354665e-7
+ ute = 2.85389809823818 lute = -8.70496079828483e-06 wute = -1.5702318701954e-06 pute = 3.78477809853975e-12
+ ua1 = 3.59568907585836e-09 lua1 = -7.04314983276821e-15 wua1 = -1.70247283463846e-15 pua1 = 3.30846469737417e-21
+ ub1 = -1.07554373303467e-18 lub1 = 1.70599534714458e-24 wub1 = 8.43397629167203e-25 pub1 = -8.01378007557458e-31
+ uc1 = -7.79450885908582e-10 luc1 = 1.66231885335503e-15 wuc1 = 3.86726099301673e-16 puc1 = -7.80861315276469e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.103 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 4.2e-07 wmax = 5.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.004443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.05323975815205+0*(0.005856/sqrt(l*w*mult))} lvth0 = 1.34039888794637e-07 wvth0 = 2.24041479748154e-09 pvth0 = -4.26225338843454e-14
+ k1 = 0.296664741042692 lk1 = 3.2976000709774e-07 wk1 = 7.04525785461585e-08 pk1 = -1.55575037829876e-13
+ k2 = 0.0594185680367042 lk2 = -1.10853872263255e-07 wk2 = -2.42379048152482e-08 pk2 = 5.32536871826916e-14
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -736385.081480147 lvsat = 1.40915481314434 wvsat = 0.369246368603152 pvsat = -6.62217143378412e-7
+ ua = -1.11166001428523e-10 lua = -1.97452069416628e-16 wua = -7.65684915258714e-17 pua = -3.37821020035555e-22
+ ub = 1.62103739275318e-18 lub = -1.29905361838012e-24 wub = -2.40452539420981e-25 pub = 7.96223089344296e-31
+ uc = -1.09088769677893e-10 luc = 1.53319609046787e-16 wuc = 9.41781431757296e-19 puc = -4.28188558585991e-23
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0142690965237155 lu0 = -5.70268546602359e-09 wu0 = -1.09833920409283e-10 pu0 = 2.04680848312011e-16
+ a0 = -0.657346400237806 la0 = 2.92102632182118e-06 wa0 = 1.05551235983987e-06 pa0 = -1.68108628811733e-12
+ keta = -0.0962974342888177 lketa = 1.26798662456746e-07 wketa = 5.10577931087838e-08 pketa = -6.90415186675651e-14
+ a1 = 0.0
+ a2 = 2.63306682296493 la2 = -3.65392175475526e-06 wa2 = -8.61068842166555e-07 pa2 = 1.71640124370659e-12
+ ags = 2.81114770247909 lags = -3.00317168385118e-06 wags = -1.27277614170947e-06 pags = 1.65982050580812e-12
+ b0 = -5.25142763609967e-07 lb0 = 1.04042517017215e-12 wb0 = 2.18024251526664e-13 pb0 = -4.54078240025689e-19
+ b1 = 1.09739058232129e-09 lb1 = -4.77784774770859e-14 wb1 = 1.03353572269177e-15 pb1 = 2.57119051808802e-20
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.532927081890699+0*(0.0/sqrt(l*w*mult))} lvoff = 7.3085599170493e-07 wvoff = 1.08323637791168e-07 pvoff = -3.83020344197045e-13
+ nfactor = {-9.72207363067639+0*(0.1/sqrt(l*w*mult))} lnfactor = 2.32551616713443e-05 wnfactor = 5.62571958286487e-06 pnfactor = -1.08880680984084e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 2.80670076923077e-05 wcit = -1.08355469408015e-11
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = -0.485738951 leta0 = 9.69238578108438e-07 weta0 = 8.97490964620035e-23 peta0 = 1.73549399148623e-29
+ etab = -0.133215546236516 letab = 2.64546941504003e-07 wetab = 1.77595448696852e-07 petab = -3.54007756514485e-13
+ dsub = 0.26
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -2.36833106801906 lpclm = 3.19218178952168e-06 wpclm = 1.37585757763034e-06 ppclm = -1.46627579749537e-12
+ pdiblc1 = 0.375532411367276 lpdiblc1 = 2.8838794189978e-08 wpdiblc1 = 8.37391601679077e-09 ppdiblc1 = -1.66920450050777e-14
+ pdiblc2 = -0.00694737337995754 lpdiblc2 = 7.32822531850026e-09 wpdiblc2 = 4.2558372800508e-09 ppdiblc2 = -4.2274848920911e-15
+ pdiblcb = 1.61421371917477 lpdiblcb = -1.82696087737763e-06 wpdiblcb = -8.63956298715339e-07 ppdiblcb = 8.58200621853297e-13
+ drout = -0.293282617079853 ldrout = 1.70088066536472e-06 wdrout = 3.16124160971165e-07 pdrout = -6.3014230278194e-13
+ pscbe1 = 720796371.089311 lpscbe1 = 157.879603245575 wpscbe1 = 48.2188649321583 ppscbe1 = -9.6116495786139e-5
+ pscbe2 = 1.07385106109966e-08 lpscbe2 = -1.86000686110179e-15 wpscbe2 = -4.15701856385516e-16 ppscbe2 = 4.97246589505542e-22
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -6.51708125521674e-11 lalpha0 = 1.64070444598945e-16 walpha0 = -1.60477968823172e-17 palpha0 = 1.59408864594873e-23
+ alpha1 = -9.93384736988146e-11 lalpha1 = 1.98010480787033e-16 walpha1 = 2.19543356333498e-21 palpha1 = -2.18080758493604e-27
+ beta0 = -202.001639105538 lbeta0 = 0.000214163831202762 wbeta0 = 0.000120014348768806 pbeta0 = -1.22595061619543e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 4.93120100905639e-10 lagidl = -2.85212285766503e-15 wagidl = -2.5029874205964e-16 pagidl = 2.04070877929026e-21
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.612971427072123 lkt1 = -8.12183203712924e-09 wkt1 = 8.99248466810301e-08 pkt1 = -2.82589588064781e-14
+ kt2 = -0.0823008217827673 lkt2 = 3.35144258515645e-08 wkt2 = 1.61961184889002e-08 pkt2 = -2.27358070273956e-14
+ at = -285745.954619788 lat = 0.402584132230619 wat = 0.175741811221126 pat = -2.02413490851081e-7
+ ute = -4.80412804441945 lute = 6.56007371686806e-06 wute = 1.8345313272009e-06 pute = -3.00206576383179e-12
+ ua1 = -4.92774614406621e-09 lua1 = 9.94693748164577e-15 wua1 = 2.34711129722896e-15 pua1 = -4.76372523687416e-21
+ ub1 = 4.74651126714728e-18 lub1 = -9.8993281228081e-24 wub1 = -1.93965598315137e-24 pub1 = 4.74618851391443e-30
+ uc1 = 2.19826576922288e-10 luc1 = -3.29578885849329e-16 wuc1 = -7.51402056895185e-17 puc1 = 1.39794341382063e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.104 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 4.2e-07 wmax = 5.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.004443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.929538946383667+0*(0.005856/sqrt(l*w*mult))} lvth0 = 1.11631718342592e-08 wvth0 = -5.4964212802604e-08 pvth0 = 1.42009964866698e-14
+ k1 = 0.630546320307838 lk1 = -1.89725308634148e-09 wk1 = -1.17911411146093e-07 pk1 = 3.15340709630451e-14
+ k2 = -0.0744147757271736 lk2 = 2.20878737644675e-08 wk2 = 4.78142506842441e-08 pk2 = -1.83184568568631e-14
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1224630.18569422 lvsat = -0.538796170320113 wvsat = -0.565442052593856 pvsat = 2.66244383556583e-7
+ ua = 1.7437277263007e-09 lua = -2.03998849513171e-15 wua = -1.17764438945664e-15 pua = 7.55919510263201e-22
+ ub = -1.31968190557306e-18 lub = 1.62207460798067e-24 wub = 1.17588856953012e-24 pub = -6.10682355138975e-31
+ uc = 7.04290413656642e-11 luc = -2.50022543395987e-17 wuc = -6.43353278308326e-17 puc = 2.20233773020835e-23
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.015596832330387 lu0 = -7.02157589675105e-09 wu0 = -2.18570454592174e-09 pu0 = 2.26672202371729e-15
+ a0 = 3.88213283914244 la0 = -1.58821090686632e-06 wa0 = -1.52640052182606e-06 pa0 = 8.83625889930946e-13
+ keta = -0.0136291570794238 lketa = 4.46811213101213e-08 wketa = 1.43239539183507e-08 pketa = -3.25524003138186e-14
+ a1 = 0.0
+ a2 = -2.86613364592984 la2 = 1.80864304061574e-06 wa2 = 1.72213768433311e-06 pa2 = -8.49595960913526e-13
+ ags = 0.205452758186985 lags = -4.14835879277947e-07 wags = -7.81936461609589e-08 pags = 4.73196318844951e-13
+ b0 = 1.05776915715599e-06 lb0 = -5.31941391377661e-13 wb0 = -5.01565532153337e-13 pb0 = 2.60717636515436e-19
+ b1 = -1.76668707943005e-07 lb1 = 1.28803343299865e-13 wb1 = 9.36586059413534e-14 pb1 = -6.62960968199847e-20
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {0.543928462211681+0*(0.0/sqrt(l*w*mult))} lvoff = -3.3882554076264e-07 wvoff = -4.29971325786959e-07 pvoff = 1.51688498333726e-13
+ nfactor = {26.6788220307582+0*(0.1/sqrt(l*w*mult))} lnfactor = -1.29032312231938e-05 wnfactor = -1.16780628019204e-05 pnfactor = 6.3004364881294e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 4.58932905741231e-05 lcit = -1.77075241852567e-11 wcit = -2.15267210541638e-11 pcit = 1.06199495114191e-17
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.49
+ etab = 0.264455062624831 letab = -1.30474385761109e-07 wetab = -3.55197579377524e-07 petab = 1.75235804406859e-13
+ dsub = 0.362722469101819 ldsub = -1.02038132012663e-07 wdsub = -8.38850903282632e-08 pdsub = 8.33262478564963e-14
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.14709555320472 lpclm = -2.9982505955151e-07 wpclm = -2.53232200968339e-07 ppclm = 1.5196098499829e-13
+ pdiblc1 = 1.16248500716365 lpdiblc1 = -7.52871123413203e-07 wpdiblc1 = -3.47988759059294e-07 ppdiblc1 = 3.3729654192965e-13
+ pdiblc2 = 0.00312009841161141 lpdiblc2 = -2.67217697599325e-09 wpdiblc2 = -1.91307069884681e-09 ppdiblc2 = 1.90032582185109e-15
+ pdiblcb = 0.488051315272615 lpdiblcb = -7.08300967410269e-07 wpdiblcb = -4.27646964534492e-07 ppdiblcb = 4.24797980456763e-13
+ drout = 2.07718519040376 ldrout = -6.53795085585443e-07 wdrout = -6.81629508084012e-07 pdrout = 3.60964331329991e-13
+ pscbe1 = 958407257.821378 lpscbe1 = -78.1483197590833 wpscbe1 = -96.4377298643171 ppscbe1 = 4.75763967758022e-5
+ pscbe2 = 4.61851862848446e-08 lpscbe2 = -3.70705367816107e-14 wpscbe2 = -1.75585125069213e-14 ppscbe2 = 1.75258518354874e-20
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 18.9476478061772 lbeta0 = -5.31349155954798e-06 wbeta0 = -7.28230508206667e-06 pbeta0 = 3.85354192337513e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -3.8544990789564e-09 lagidl = 1.46653248322078e-15 wagidl = 2.86797340045364e-15 pagidl = -1.05678943420959e-21
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.731406532524195 lkt1 = 1.09524258742421e-07 wkt1 = 1.22133617091925e-07 pkt1 = -6.0253154388896e-14
+ kt2 = -0.100048195293156 lkt2 = 5.11435663596272e-08 wkt2 = 3.3583486092534e-08 pkt2 = -4.00073399880541e-14
+ at = 125974.305421817 lat = -0.00639324743858949 wat = -0.0278044992997943 pat = -2.23205850851177e-10
+ ute = 3.48358389471905 lute = -1.6724254853319e-06 wute = -2.24969242817295e-06 pute = 1.05494889288376e-12
+ ua1 = 1.00853785738006e-08 lua1 = -4.96616979935064e-15 wua1 = -5.03818960486036e-15 pua1 = 2.57237479060544e-21
+ ub1 = -1.08912684714139e-17 lub1 = 5.63427272713478e-24 wub1 = 5.66995620747082e-24 pub1 = -2.81272844029384e-30
+ uc1 = -2.46429547484996e-10 luc1 = 1.33571040257153e-16 wuc1 = 1.30309439485697e-16 puc1 = -6.42865982569946e-23
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.105 pmos
* DC IV MOS Parameters
+ lmin = 2.5e-07 lmax = 5e-07 wmin = 4.2e-07 wmax = 5.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.006443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.853457644131067+0*(0.007356/sqrt(l*w*mult))} lvth0 = -2.63706256564339e-08 wvth0 = -5.1659753315767e-08 pvth0 = 1.25707810523522e-14
+ k1 = 0.671917546540906 lk1 = -2.23072510937112e-08 wk1 = -1.06544435155784e-07 pk1 = 2.59263097619382e-14
+ k2 = -0.0443411185594837 lk2 = 7.25139588467364e-09 wk2 = 2.10805197888021e-08 pk2 = -5.12969152436754e-15
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 152097.532347528 lvsat = -0.00967505618336287 wvsat = -0.0508386711438604 pvsat = 1.23709805588047e-8
+ ua = -3.21176728642792e-09 lua = 4.04745503457798e-16 wua = 6.9977112982976e-16 pua = -1.70280907190514e-22
+ ub = 2.24513110982347e-18 lub = -1.36583115409023e-25 wub = -1.22287360096497e-25 pub = 2.97571616311615e-32
+ uc = 3.89183171258982e-11 luc = -9.45681666460102e-18 wuc = -3.88627386372953e-17 puc = 9.45678109452218e-24
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = -0.00270245356241038 lu0 = 2.00615720702982e-09 wu0 = 4.75372365776541e-09 pu0 = -1.15676160743332e-15
+ a0 = 0.517502082202142 la0 = 7.16893015010951e-08 wa0 = 5.22378037177278e-07 pa0 = -1.27114426810645e-13
+ keta = 0.161533335343541 lketa = -4.17331923768395e-08 wketa = -1.01943398142589e-07 pketa = 2.48067026172214e-14
+ a1 = 0.0
+ a2 = 1.06891451743248 la2 = -1.32665750201105e-7
+ ags = -1.66447624457111 lags = 5.07671155084724e-07 wags = 1.73848168734078e-06 pags = -4.23038656834131e-13
+ b0 = -4.04146836985534e-08 lb0 = 9.83442830183858e-15 wb0 = 5.31052000558932e-14 pb0 = -1.29225131712009e-20
+ b1 = 1.66583825042715e-07 lb1 = -4.05361748182441e-14 wb1 = -8.03629899283572e-14 pb1 = 1.95553692431866e-20
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {0.128997699621305+0*(0.0/sqrt(l*w*mult))} lvoff = -1.34124428207829e-07 wvoff = -2.41730782349445e-07 pvoff = 5.88222851153493e-14
+ nfactor = {-1.90807716553442+0*(0.1/sqrt(l*w*mult))} lnfactor = 1.19977245250681e-06 wnfactor = 2.15681736622238e-06 pnfactor = -5.24835624261821e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.49
+ etab = 2.62181963977308e-05 letab = -2.1588508475031e-11 wetab = 1.33639676417029e-11 petab = -3.2519611579967e-18
+ dsub = -0.30363875647572 ldsub = 2.26703182291309e-07 wdsub = 1.67770180656526e-07 pdsub = -4.08248602205979e-14
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.444148646507052 lpclm = 4.69653615049074e-08 wpclm = 1.08127669747885e-07 ppclm = -2.63115709011107e-14
+ pdiblc1 = -1.16713263793553 lpdiblc1 = 3.96417786384735e-07 wpdiblc1 = 6.62481854051425e-07 ppdiblc1 = -1.61207009401166e-13
+ pdiblc2 = -0.0153041644819908 lpdiblc2 = 6.41721203141068e-09 wpdiblc2 = 3.82614139769362e-09 ppdiblc2 = -9.31045595431972e-16
+ pdiblcb = -1.65110263054523 lpdiblcb = 3.47024961911615e-07 wpdiblcb = 8.55293929068984e-07 ppdiblcb = -2.08125514111788e-13
+ drout = 1.0636610152262 ldrout = -1.53785096051692e-07 wdrout = 9.87623722833648e-08 pdrout = -2.40326381466894e-14
+ pscbe1 = 800069244.26128 lpscbe1 = -0.034160825371373
+ pscbe2 = -6.61067699640808e-08 lpscbe2 = 1.83273523303217e-14 wpscbe2 = 3.54542815693916e-14 ppscbe2 = -8.62737396853262e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 7.09089376038267 lbeta0 = 5.358957678962e-07 wbeta0 = 1.04361639519408e-06 pbeta0 = -2.53951526373735e-13
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -1.83748873357367e-09 lagidl = 4.71464633450349e-16 wagidl = 1.43236330889361e-15 pagidl = -3.48548422859554e-22
+ bgidl = 730034204.0064 lbgidl = 133.184385863891
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.506801150159999 lkt1 = -1.28211138236582e-9
+ kt2 = 0.0242671675443682 lkt2 = -1.01859261119115e-08 wkt2 = -9.3757320504542e-08 pkt2 = 2.28147188569342e-14
+ at = 158236.242086396 lat = -0.0223092867488195 wat = -0.0557608877056524 pat = 1.3568742892518e-8
+ ute = 0.364968229524015 lute = -1.33893870295915e-07 wute = -2.19639480984915e-07 pute = 5.34466320239072e-14
+ ua1 = -3.54490332115945e-10 lua1 = 1.8421424695643e-16 wua1 = 3.47377629291368e-16 pua1 = -8.45301775565029e-23
+ ub1 = 6.17482959937584e-19 lub1 = -4.34316865052916e-26 wub1 = -6.20943392504082e-26 pub1 = 1.51099123245158e-32
+ uc1 = 4.743483235632e-11 luc1 = -1.14034251650022e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.24e-6
+ sbref = 1.24e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.106 pmos
* DC IV MOS Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 4.2e-07 wmax = 5.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.006443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.772463663771427+0*(0.007356/sqrt(l*w*mult))} lvth0 = -4.60795388491878e-8
+ k1 = -0.415479539169429 lk1 = 2.4229778094887e-7
+ k2 = 0.438589349394085 lk2 = -1.10263938326212e-07 pk2 = -2.20881053461883e-29
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 92623.7868717143 lvsat = 0.00479716609323078
+ ua = -1.55915274021429e-09 lua = 2.60158501126512e-18
+ ub = 9.27892318000016e-20 lub = 3.87163452505452e-25
+ uc = 6.09622494694279e-15 luc = 1.20053449946548e-20
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0028191509837143 lu0 = 6.62540999984935e-10
+ a0 = -0.39776447742857 la0 = 2.94408435588514e-7
+ keta = -0.184161871607297 lketa = 4.23875878921637e-08 wketa = 1.32348898008484e-23
+ a1 = 0.0
+ a2 = 0.164955374458 la2 = 8.73018597320193e-8
+ ags = -1.62902379023886 lags = 4.99044225752423e-7
+ b0 = 1.23812857142857e-09 lb0 = -3.01283730314285e-16
+ b1 = -1.86798933828571e-10 lb1 = 4.54552789599769e-17
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.403685441391143+0*(0.0/sqrt(l*w*mult))} lvoff = -4.50237804014202e-9
+ nfactor = {-5.59783716277429+0*(0.1/sqrt(l*w*mult))} lnfactor = 2.09763127071517e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 1.39713389074943 leta0 = -2.20740146707184e-07 peta0 = 1.0097419586829e-28
+ etab = 0.244655617911143 letab = -5.95492173762617e-08 wetab = 2.98818996284781e-23 petab = 3.10613981430773e-30
+ dsub = 1.53653693089571 ldsub = -2.21081489122281e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.664807054980857 lpclm = -6.72921429629188e-9
+ pdiblc1 = 1.18699067550629 lpdiblc1 = -1.76429872461569e-07 wpdiblc1 = -4.2351647362715e-22
+ pdiblc2 = 0.0300992129326343 lpdiblc2 = -4.63115502190936e-9
+ pdiblcb = -0.782143533009561 lpdiblcb = 1.3557419303548e-7
+ drout = -0.975627884693999 ldrout = 3.42451386277088e-7
+ pscbe1 = 799752699.066858 lpscbe1 = 0.0428666491488912
+ pscbe2 = 2.95389305828885e-08 lpscbe2 = -4.94688114937674e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 11.56376242988 lbeta0 = -5.52523148401942e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -1.10815918728486e-08 lagidl = 2.72090620315523e-15 wagidl = -2.95822839457879e-31 pagidl = -1.17549435082229e-37
+ bgidl = 1964163557.12 lbgidl = -167.126182664067
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.238369297999999 lkt1 = -6.66017814232761e-8
+ kt2 = 0.235996541485714 lkt2 = -6.17077285080507e-08 wkt2 = -2.64697796016969e-23 pkt2 = 3.15544362088405e-30
+ at = -4339.24200000009 lat = 0.017251506397796
+ ute = -0.316907829714286 lute = 3.20324862070148e-8
+ ua1 = 9.89437705428572e-10 lua1 = -1.42814513843578e-16 wua1 = 3.94430452610506e-31
+ ub1 = 6.03324424e-19 lub1 = -3.99863766873121e-26
+ uc1 = -5.82329727011428e-11 luc1 = 1.43095671820707e-17 wuc1 = -1.23259516440783e-32 puc1 = -2.57139389242375e-39
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.107 pmos
* DC IV MOS Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 4.2e-07 wmax = 5.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+0*(4.01004e-09*(0.006443/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.271654364967343+0*(0.007356/sqrt(l*w*mult))} lvth0 = -1.32888821085291e-07 wvth0 = -3.98278310386429e-07 pvth0 = 6.90367657657628e-14
+ k1 = -3.55748906215231 lk1 = 7.86927427643677e-07 wk1 = 2.03056188465519e-06 pk1 = -3.51973535962361e-13
+ k2 = 0.776126409588245 lk2 = -1.68771937266147e-07 wk2 = -4.41168841059264e-07 pk2 = 7.64713245715306e-14
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 726436.861837209 lvsat = -0.105066724695138 wvsat = -0.291535788567276 pvsat = 5.05342305186745e-8
+ ua = 3.56276519618137e-09 lua = -8.85221426247687e-16 wua = -1.77835174337371e-16 pua = 3.08255934492912e-23
+ ub = 8.79862749666121e-19 lub = 2.50733703065572e-25 wub = -3.2510133643624e-25 pub = 5.63524154551854e-32
+ uc = 8.50235402252939e-13 luc = -1.34316051721212e-19 wuc = -7.01400254704987e-19 puc = 1.21579317350053e-25
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0249695907796761 lu0 = -3.1769719333675e-09 wu0 = -6.3668616419242e-10 pu0 = 1.10361906328787e-16
+ a0 = 8.32068401515669 la0 = -1.21682998921923e-06 wa0 = -2.3328071300386e-06 pa0 = 4.04364122306631e-13
+ keta = 1.11264356092967 lketa = -1.8239807217293e-07 wketa = -3.86463345221317e-07 pketa = 6.69887833339726e-14
+ a1 = 0.0
+ a2 = -4.40683997149522 la2 = 8.7976772140886e-07 wa2 = 2.66744726566008e-06 pa2 = -4.62369974134988e-13
+ ags = -12.5265781191666 lags = 2.3880044980201e-06 wags = 6.47144011416919e-06 pags = -1.12174648650986e-12
+ b0 = -9.43786834473983e-06 lb0 = 1.63585455414051e-12 wb0 = 3.70922238735812e-12 pb0 = -6.42949190179883e-19
+ b1 = -1.58275104845512e-07 lb1 = 2.74481660490793e-14 wb1 = 2.83500848521524e-14 pb1 = -4.9141470081024e-21
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.2417827539422+0*(0.0/sqrt(l*w*mult))} lvoff = 1.40771733922834e-07 wvoff = 5.43094333486554e-07 pvoff = -9.41388855778923e-14
+ nfactor = {9.86831059126987+0*(0.1/sqrt(l*w*mult))} lnfactor = -5.83239848675335e-07 wnfactor = -2.25723831182213e-07 pnfactor = 3.91265174494643e-14
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = -1.9160829999519 leta0 = 3.53566242693203e-07 weta0 = 1.06293107742129e-06 peta0 = -1.84246347098052e-13
+ etab = -0.883950891803182 letab = 1.360811778046e-07 wetab = 2.51387450396963e-07 petab = -4.35749978769088e-14
+ dsub = 0.266362313510667 ldsub = -9.11961293991947e-10
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 3.60108054627701 lpclm = -5.15696988730585e-07 wpclm = -1.76002110450694e-06 ppclm = 3.05078538213025e-13
+ pdiblc1 = 2.54722785653482 lpdiblc1 = -4.12210664946693e-07 wpdiblc1 = -1.45126962854731e-06 ppdiblc1 = 2.51560174873133e-13
+ pdiblc2 = 0.0582974018945875 lpdiblc2 = -9.51897270019641e-09 wpdiblc2 = -3.36595131794213e-08 ppdiblc2 = 5.83447269549454e-15
+ pdiblcb = 1.65062695831742 lpdiblcb = -2.86117378390157e-07 wpdiblcb = -7.75056069871773e-07 ppdiblcb = 1.34346669039433e-13
+ drout = -0.559222936309904 ldrout = 2.70272585334086e-07 wdrout = 9.35131794112962e-07 pdrout = -1.62093874927952e-13
+ pscbe1 = 748810658.381924 lpscbe1 = 8.87305809739428 wpscbe1 = 30.7004083585762 ppscbe1 = -5.32154738405884e-6
+ pscbe2 = -6.16991658561486e-08 lpscbe2 = 1.08681480111731e-14 wpscbe2 = 1.35276716553977e-14 ppscbe2 = -2.34485954940332e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 28.0186167079081 lbeta0 = -3.40477467924677e-06 wbeta0 = -1.00152266064487e-05 pbeta0 = 1.73601934950861e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 2.56215189917322e-08 lagidl = -3.64113762788948e-15 wagidl = -3.70937252476877e-15 pagidl = 6.4297521469837e-22
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.186819280934522 lkt1 = -7.55373582813718e-08 wkt1 = -2.04704593691399e-07 pkt1 = 3.54830848612796e-14
+ kt2 = -0.12
+ at = 367446.271380506 lat = -0.0471930509205542 wat = -0.0586053616739162 pat = 1.01585361818333e-8
+ ute = -3.56208572623696 lute = 5.94545132434462e-07 wute = 1.67853625105275e-06 pute = -2.90954116684981e-13
+ ua1 = -1.25921172055398e-10 lua1 = 5.05195632617386e-17 wua1 = 2.15887242208684e-16 pua1 = -3.74214627899689e-23
+ ub1 = 3.7264e-19
+ uc1 = 2.53798686275156e-10 luc1 = -3.97773765215631e-17 wuc1 = -1.38499172747403e-16 puc1 = 2.40071696056894e-23
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.29e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+2.0e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+4.5e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+2.5e-7}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.5}
+ steta0 = 0.0
+ tku0 = 0.0
.ends sky130_fd_pr__pfet_01v8
