* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
.subckt  sky130_fd_pr__pfet_g5v0d10v5 d g s b
+ 
.param  l = 1 w = 1 ad = 0 as = 0 pd = 0 ps = 0 nrd = 0 nrs = 0 sa = 0 sb = 0 sd = 0 mult = 1 nf = 1.0
msky130_fd_pr__pfet_g5v0d10v5 d g s b sky130_fd_pr__pfet_g5v0d10v5__model l = {l} w = {w} ad = {ad} as = {as} pd = {pd} ps = {ps} nrd = {nrd} nrs = {nrs} sa = {sa} sb = {sb} sd = {sd} nf = {nf}
.model sky130_fd_pr__pfet_g5v0d10v5__model.0 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 2.0e-05 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.979018+0*(0.0/sqrt(l*w*mult))}
+ k1 = 0.59521
+ k2 = 0.0218501
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200000.0
+ ua = 2.70482362e-9
+ ub = -1.668e-20
+ uc = -3.9972e-11
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0213783
+ a0 = 0.8929174
+ keta = -0.0079259
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.145547
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.093204657+0*(0.009/sqrt(l*w*mult))}
+ nfactor = {1.76562+0*(0.02/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.0800000000000101
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.08353125
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0029407877
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 333712830.0
+ pscbe2 = 1.5000958e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 5.0667189e-5
+ alpha1 = 0.0
+ beta0 = 38.266046
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 7.3657e-9
+ bgidl = 1704700000.0
+ cgidl = 700.0
+ egidl = 0.69350825
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.57573
+ kt2 = -0.019032
+ at = 430000.0
+ ute = -1.3864
+ ua1 = 7.0656e-10
+ ub1 = -3.145e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.1 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 2.0e-05 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.979018+0*(0.0/sqrt(l*w*mult))}
+ k1 = 0.59521
+ k2 = 0.0218501
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200000.0
+ ua = 2.70482362e-9
+ ub = -1.668e-20
+ uc = -3.9972e-11
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0213783
+ a0 = 0.8929174
+ keta = -0.0079259
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.145547
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.093204657+0*(0.009/sqrt(l*w*mult))}
+ nfactor = {1.76562+0*(0.02/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.0800000000000101
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.08353125
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0029407877
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 333712830.0
+ pscbe2 = 1.5000958e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 5.0667189e-5
+ alpha1 = 0.0
+ beta0 = 38.266046
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 7.3657e-9
+ bgidl = 1704700000.0
+ cgidl = 700.0
+ egidl = 0.69350825
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.57573
+ kt2 = -0.019032
+ at = 430000.0
+ ute = -1.3864
+ ua1 = 7.0656e-10
+ ub1 = -3.145e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.2 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 2.0e-05 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.98502420227+0*(0.0/sqrt(l*w*mult))} lvth0 = 4.7358874867938e-8
+ k1 = 0.6040969260625 lk1 = -7.0073367568183e-8
+ k2 = 0.019548143337625 lk2 = 1.81509167730436e-8
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 297115.1625125 lvsat = -0.76575257083525
+ ua = 2.45140613429905e-09 lua = 1.99819560766456e-15
+ ub = 2.39982194675e-19 lub = -2.0237801217014e-24 wub = -9.18354961579912e-41 pub = -3.50324616081204e-45
+ uc = -5.150363640875e-11 luc = 9.09268954248118e-17
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.02071299460625 lu0 = 5.2459297031918e-9
+ a0 = 0.912995345534625 la0 = -1.58314500150792e-7
+ keta = -0.004975149172625 lketa = -2.32666555200977e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.1193446512225 lags = 2.06605389098844e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0947667260771125+0*(0.009/sqrt(l*w*mult))} lvoff = 1.23169068626866e-8
+ nfactor = {1.7731568903+0*(0.02/sqrt(l*w*mult))} lnfactor = -5.94283423310471e-8
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.0800000000000101
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.643778489125225 lpclm = 5.7348336564537e-06 wpclm = -1.6940658945086e-21 ppclm = 6.46234853557053e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00454411319014038 lpdiblc2 = -1.26422134731294e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 560706123.996462 lpscbe1 = -1789.84098819564
+ pscbe2 = -1.51292780647975e-08 lpscbe2 = 2.37576760719748e-13
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 7.7982685969875e-05 lalpha0 = -2.1538255702998e-10
+ alpha1 = 0.0
+ beta0 = 39.1348639430788 lbeta0 = -6.85062513708622e-06 wbeta0 = 2.16840434497101e-19
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 6.543926432625e-09 lagidl = 6.47968046988403e-15
+ bgidl = 1479758789.5 lbgidl = 1773.66032008645
+ cgidl = 931.1572025 lcgidl = -0.00182267338592649
+ egidl = 1.20611845100666 legidl = -4.04192887188653e-6
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.5851802503375 lkt1 = 7.45151766599359e-8
+ kt2 = -0.019032
+ at = 671539.8516375 lat = -1.90454052246243
+ ute = -1.221579087125 lute = -1.29961207391481e-6
+ ua1 = 1.37134480442e-09 lua1 = -5.24182485892768e-15
+ ub1 = -2.61372693375e-18 lub1 = -4.18908547101592e-24
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.3 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 2.0e-05 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.9582756181165+0*(0.0/sqrt(l*w*mult))} lvth0 = -5.65592408254869e-8
+ k1 = 0.6023840567 lk1 = -6.34188786592167e-8
+ k2 = 0.02423914419975 lk2 = -7.35981213077727e-11
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 84741.5405 lvsat = 0.0593178888152026
+ ua = 3.31429591882863e-09 lua = -1.35412689078391e-15
+ ub = -1.22040265805e-18 lub = 3.64980772921096e-24 wub = -2.93873587705572e-39
+ uc = -5.45822372525e-11 luc = 1.02887244309776e-16
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0211909620139 lu0 = 3.38902871430858e-9
+ a0 = 0.82381514871175 la0 = 1.88150118605095e-7
+ keta = -0.00516198539 lketa = -2.2540797749777e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.1427222865525 lags = 1.1578339272997e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0644364973897325+0*(0.009/sqrt(l*w*mult))} lvoff = -1.05515879936641e-7
+ nfactor = {2.19899029989+0*(0.02/sqrt(l*w*mult))} lnfactor = -1.71378900942115e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.0198686595000102 leta0 = 2.33609957185798e-7
+ etab = -0.12173557277 letab = 2.00992441533586e-7
+ dsub = 0.811505457875 ldsub = -9.77097446317086e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.04601663892438 lpclm = -8.30011967043352e-7
+ pdiblc1 = 0.5791285228315 lpdiblc1 = -7.34763365557763e-7
+ pdiblc2 = -0.00110255629368 lpdiblc2 = 9.29506923816533e-09 ppdiblc2 = -2.52435489670724e-29
+ pdiblcb = 0.1634995 lpdiblcb = -7.323196150025e-07 wpdiblcb = 4.2351647362715e-22 ppdiblcb = -1.21169035041947e-27
+ drout = 0.1453011 ldrout = 1.6111031530055e-6
+ pscbe1 = -152915980.78355 lpscbe1 = 982.577320764188
+ pscbe2 = 7.56929177375625e-08 lpscbe2 = -1.15267015861442e-13
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 4.37897997750275e-05 lalpha0 = -8.2543365127428e-11
+ alpha1 = -9.424975e-11 lalpha1 = 3.6615980750125e-16
+ beta0 = 69.7665703037275 lbeta0 = -0.000125854651189675
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 9.1846459195e-09 lagidl = -3.7795015330279e-15
+ bgidl = 2611316709.5 lbgidl = -2622.43654132395
+ cgidl = 455.826641375 lcgidl = 2.39834673913318e-5
+ egidl = -1.56307736015895 legidl = 6.71638300851282e-06 wegidl = 3.3881317890172e-21 pegidl = 6.46234853557053e-27
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.5669424975 lkt1 = 3.6615980750127e-9
+ kt2 = -0.019032
+ at = 210065.598725 lat = -0.111715357268631
+ ute = -1.70322385975 lute = 5.71575459509452e-7
+ ua1 = -4.7771419424e-10 lua1 = 1.94176010557143e-15 wua1 = 7.88860905221012e-31 pua1 = 1.50463276905253e-36
+ ub1 = -3.71961517675e-18 lub1 = 1.07284823597865e-25
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.4 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 2.0e-05 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.0103795446465+0*(0.0/sqrt(l*w*mult))} lvth0 = 4.1656400163929e-8
+ k1 = 0.55931480325 lk1 = 1.77664487477661e-8
+ k2 = 0.0189737620275 lk2 = 9.85162094647264e-9
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 176673.743395 lvsat = -0.113973853980858
+ ua = 3.433765183409e-09 lua = -1.5793258571716e-15
+ ub = 6.855908709e-19 lub = 5.70194571078546e-26
+ uc = 5.181291727e-13 luc = -9.76670899893637e-19
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0261944534892 lu0 = -6.04252769917455e-9
+ a0 = 0.9866834812625 la0 = -1.18855873911406e-7
+ keta = 0.04266318224 lketa = -1.12690999606489e-07 pketa = 1.0097419586829e-28
+ a1 = 0.0
+ a2 = 0.5
+ ags = -0.3008568383605 lags = 9.51927825295351e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.158164876157715+0*(0.009/sqrt(l*w*mult))} lvoff = 7.1161645399112e-8
+ nfactor = {1.03928807542+0*(0.02/sqrt(l*w*mult))} lnfactor = 4.72243885193677e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.4424975e-05 lcit = -8.341055750125e-12
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.271036933858215 leta0 = -2.39840984138047e-7
+ etab = -0.02847850446 letab = 2.52033340545777e-8
+ dsub = 0.0710074050500002 ldsub = 4.18737680767775e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.0769866827459003 lpclm = 9.96604655203293e-7
+ pdiblc1 = 0.0033121379690001 lpdiblc1 = 3.50647640826125e-7
+ pdiblc2 = 0.0058837902087835 lpdiblc2 = -3.87415898724585e-9
+ pdiblcb = -0.401999 lpdiblcb = 3.33642230005e-7
+ drout = 1.52153692559705 ldrout = -9.83094497065811e-7
+ pscbe1 = 429292893.4686 lpscbe1 = -114.883496156744
+ pscbe2 = 1.453303481712e-08 lpscbe2 = 1.9057644177885e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -6.0014119919695e-05 lalpha0 = 1.13126504477525e-10 walpha0 = -9.02811862980187e-26 palpha0 = -1.33339051360666e-31
+ alpha1 = 1.884995e-10 lalpha1 = -1.668211150025e-16
+ beta0 = -38.730102860375 lbeta0 = 7.86610352412926e-05 wbeta0 = -5.42101086242752e-20
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 3.931314352e-09 lagidl = 6.12300220505176e-15
+ bgidl = 865040006.000001 lbgidl = 669.28631339003
+ cgidl = 440.29210965 lcgidl = 5.32659820202982e-5
+ egidl = 3.0805973382958 legidl = -2.03692057970089e-6
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.501988356 lkt1 = -1.1877663388178e-7
+ kt2 = -0.019032
+ at = 257884.395 lat = -0.201853549153025
+ ute = -1.2168945345 lute = -3.45152886940173e-7
+ ua1 = 6.697326371e-10 lua1 = -2.21171434270314e-16
+ ub1 = -3.5355262185e-18 lub1 = -2.39721942258593e-25
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.81e-6
+ sbref = 2.81e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.5 pmos
* DC IV MOS Parameters
+ lmin = 8.0e-07 lmax = 1e-06 wmin = 2.0e-05 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.0629626301025+0*(0.0/sqrt(l*w*mult))} lvth0 = 8.81921678770623e-8
+ k1 = 0.589870423499999 lk1 = -9.27512239538251e-9
+ k2 = 0.0153723850424999 lk2 = 1.30388215713127e-8
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 6575.92405749997 lvsat = 0.0365618656437328
+ ua = -7.372924266755e-10 lua = 2.11203927246513e-15
+ ub = 4.0360095145e-18 lub = -2.90808429038493e-24
+ uc = 5.8546574915e-12 luc = -5.69947177939004e-18 puc = -1.17549435082229e-38
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.02041063238 lu0 = -9.23874936638109e-10
+ a0 = 0.8827697056925 la0 = -2.68927021008339e-8
+ keta = -0.15139736295 lketa = 5.90516125839353e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.9585371661525 lags = -1.62629571728632e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0946561577386999+0*(0.009/sqrt(l*w*mult))} lvoff = 1.49567471418758e-8
+ nfactor = {0.847250546749999+0*(0.02/sqrt(l*w*mult))} lnfactor = 6.42196137878983e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -1.2124875e-05 lcit = 1.5155428750625e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -6.82344178649e-05 leta0 = 8.57342604422856e-11
+ etab = 0.00072873193075 letab = -6.44924115054096e-10
+ dsub = 1.4666427665 ldsub = -8.16392635938667e-07 wdsub = -6.7762635780344e-21
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.99390052644125 lpclm = -6.99854511897874e-7
+ pdiblc1 = 0.20282696902275 lpdiblc1 = 1.74078012917712e-7
+ pdiblc2 = -0.0324173066339675 lpdiblc2 = 3.00221202131046e-08 wpdiblc2 = 2.64697796016969e-23
+ pdiblcb = -0.025
+ drout = 0.3384020931485 ldrout = 6.39739139769935e-8
+ pscbe1 = -44797159.5075004 lpscbe1 = 304.68383027684
+ pscbe2 = 1.815406017615e-08 lpscbe2 = -3.18553169343687e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.00024102438742525 lalpha0 = -1.53291069330214e-10
+ alpha1 = 0.0
+ beta0 = 66.614022720125 lbeta0 = -1.4567989176822e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 9.10326274999998e-09 lagidl = 1.54585373256375e-15
+ bgidl = 984254649.999999 lbgidl = 563.781949523251
+ cgidl = 433.624488 lcgidl = 5.916679384244e-5
+ egidl = 1.79942371219525 legidl = -9.03088326470035e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.6111976825 lkt1 = -2.21269259759127e-8
+ kt2 = -0.019032
+ at = 46239.88 lat = -0.0145492116006
+ ute = -2.0422143225 lute = 3.85250998840888e-7
+ ua1 = -3.42631855000003e-11 lua1 = 4.01861348751572e-16
+ ub1 = -4.54448211249999e-18 lub1 = 6.53198979151934e-25
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.41e-6
+ sbref = 2.41e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.6 pmos
* DC IV MOS Parameters
+ lmin = 6e-07 lmax = 8.0e-07 wmin = 2.0e-05 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.881892254404999+0*(0.0/sqrt(l*w*mult))} lvth0 = -3.58401341238466e-8
+ k1 = 0.59352307275 lk1 = -1.17771688683862e-8
+ k2 = 0.0189560867925 lk2 = 1.05840037910715e-8
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 61502.5565075 lvsat = -0.00106260295135498
+ ua = -1.8233767778005e-09 lua = 2.85600162256401e-15
+ ub = 2.469434477865e-18 lub = -1.83498822316514e-24 wub = 2.93873587705572e-39 pub = 1.40129846432482e-45
+ uc = 2.53255847e-12 luc = -3.42385056015765e-18
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.00709052591749999 lu0 = 8.20033138964209e-9
+ a0 = 0.93451931175 la0 = -6.23409235021911e-8
+ keta = 0.011718082125 lketa = -5.26816517152144e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = -0.561400778000001 lags = 8.7852032032611e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {0.00731538466477499+0*(0.009/sqrt(l*w*mult))} lvoff = -5.48932495467926e-8
+ nfactor = {1.78668573025+0*(0.02/sqrt(l*w*mult))} lnfactor = -1.31226564259881e-9
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -0.0573036120981399 leta0 = 3.92916817945423e-08 weta0 = -6.45200877791362e-23 peta0 = -1.97215226305253e-29
+ etab = -0.00072873193075 letab = 3.53431342754096e-10
+ dsub = 0.1933921039715 ldsub = 5.57777016400423e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.25744420752125 lpclm = 4.89609384280732e-7
+ pdiblc1 = 0.18971742632875 lpdiblc1 = 1.83057984115388e-7
+ pdiblc2 = 0.02598707339889 lpdiblc2 = -9.98458808750266e-9
+ pdiblcb = -0.025
+ drout = -0.6825930358415 ldrout = 7.63350472359499e-7
+ pscbe1 = 430689610.609 lpscbe1 = -21.0222298191119
+ pscbe2 = 1.0686514267575e-08 lpscbe2 = 1.92969991620746e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -0.000115023676316125 lalpha0 = 9.06000740923091e-11 walpha0 = 2.06795153138257e-25
+ alpha1 = 0.0
+ beta0 = 27.36521542835 lbeta0 = 1.23172475740074e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 2.30942115275e-08 lagidl = -8.03787622527987e-15
+ bgidl = 2050039997.5 lbgidl = -166.275684587513
+ cgidl = 1223.24275 lcgidl = -0.00048171776753625
+ egidl = -0.212081994370001 legidl = 4.74783024998628e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.7041728745 lkt1 = 4.15606156681274e-8
+ kt2 = -0.019032
+ at = 41974.825 lat = -0.011627670250875
+ ute = -1.6071111875 lute = 8.72075268815624e-8
+ ua1 = 5.5336999e-10 lua1 = -6.64438300050192e-19
+ ub1 = -4.2982652075e-18 lub1 = 4.84541630311462e-25
+ uc1 = -2.733805074e-10 luc1 = 1.12462826666463e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.02e-6
+ sbref = 2.01e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.7 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 6e-07 wmin = 2.0e-05 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.02/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.862969830475+0*(0.0/sqrt(l*w*mult))} lvth0 = -4.50174151177776e-8
+ k1 = 0.45836144 lk1 = 5.37755472072001e-8
+ k2 = 0.0407020010000001 lk2 = 3.73441300049918e-11
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 38739.7771700001 lvsat = 0.00997723121343586
+ ua = 1.1407329461341e-08 lua = -3.56082474988843e-15
+ ub = -7.45358295523e-18 lub = 2.97762561679878e-24 wub = -2.35098870164458e-38
+ uc = -1.62221272500001e-12 luc = -1.40880730443863e-18
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.037707886955 lu0 = -6.64893562674022e-9
+ a0 = 0.214396683 la0 = 2.86914950828415e-7
+ keta = -0.13938919825 lketa = 2.06046237302588e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 1.25
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1225417579515+0*(0.009/sqrt(l*w*mult))} lvoff = 8.08681533638781e-9
+ nfactor = {1.294882352+0*(0.02/sqrt(l*w*mult))} lnfactor = 2.3720991379176e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 2.924975e-05 lcit = -9.33603250125e-12
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -0.19321058279999 leta0 = 1.05205883050086e-07 weta0 = -4.2351647362715e-22
+ etab = 0.014823462485 letab = -7.18930518791258e-9
+ dsub = 0.419003534557 ldsub = -5.36427141367724e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.998842207075001 lpclm = 1.3003506148716e-7
+ pdiblc1 = 1.618697765494 lpdiblc1 = -5.09990335478063e-7
+ pdiblc2 = 0.00770696779005001 lpdiblc2 = -1.1188282677433e-9
+ pdiblcb = -0.025
+ drout = 0.859530092143 ldrout = 1.54284659026556e-8
+ pscbe1 = 482455064.78 lpscbe1 = -46.128216264776
+ pscbe2 = 1.53528728706e-08 lpscbe2 = -3.33460674466651e-16
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -2.58245787587999e-05 lalpha0 = 4.73389577724942e-11
+ alpha1 = 0.0
+ beta0 = 45.3597691823501 lbeta0 = 3.58997897608615e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -2.1841096655e-08 lagidl = 1.37555235666917e-14
+ bgidl = 2064090365 lbgidl = -173.090042573175
+ cgidl = -2257.0677 lcgidl = 0.0012062153991615 wcgidl = 3.46944695195361e-18 pcgidl = -1.65436122510606e-24
+ egidl = 1.15799168033 legidl = -1.89695856862499e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.637729750000001 lkt1 = 9.33603250125007e-9
+ kt2 = -0.019032
+ at = 18000.0
+ ute = -1.638662255 lute = 1.02509636863725e-7
+ ua1 = 5.52e-10
+ ub1 = -7.68506304000001e-18 lub1 = 2.1271216450848e-24
+ uc1 = -4.1496e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 1.81e-6
+ sbref = 1.81e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.8 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 1.5e-05 wmax = 2.0e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.979018+0*(0.0/sqrt(l*w*mult))}
+ k1 = 0.59521
+ k2 = 0.0218501
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200000.0
+ ua = 2.70482362e-9
+ ub = -1.668e-20
+ uc = -3.9972e-11
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0213783
+ a0 = 0.8929174
+ keta = -0.0079259
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.145547
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.093204657+0*(0.009/sqrt(l*w*mult))}
+ nfactor = {1.76562+0*(0.02/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.0800000000000101
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.08353125
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0029407877
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 333712830.0
+ pscbe2 = 1.5000958e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 5.0667189e-5
+ alpha1 = 0.0
+ beta0 = 38.266046
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 7.3657e-9
+ bgidl = 1704700000.0
+ cgidl = 700.0
+ egidl = 0.69350825
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.57573
+ kt2 = -0.019032
+ at = 430000.0
+ ute = -1.3864
+ ua1 = 7.0656e-10
+ ub1 = -3.145e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.9 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 1.5e-05 wmax = 2.0e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.979018+0*(0.0/sqrt(l*w*mult))}
+ k1 = 0.59521
+ k2 = 0.0218501
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200000.0
+ ua = 2.70482362e-9
+ ub = -1.668e-20
+ uc = -3.9972e-11
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0213783
+ a0 = 0.8929174
+ keta = -0.0079259
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.145547
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.093204657+0*(0.009/sqrt(l*w*mult))}
+ nfactor = {1.76562+0*(0.02/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.0800000000000101
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.08353125
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0029407877
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 333712830.0
+ pscbe2 = 1.5000958e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 5.0667189e-5
+ alpha1 = 0.0
+ beta0 = 38.266046
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 7.3657e-9
+ bgidl = 1704700000.0
+ cgidl = 700.0
+ egidl = 0.69350825
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.57573
+ kt2 = -0.019032
+ at = 430000.0
+ ute = -1.3864
+ ua1 = 7.0656e-10
+ ub1 = -3.145e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.10 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 1.5e-05 wmax = 2.0e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.985024202269999+0*(0.0/sqrt(l*w*mult))} lvth0 = 4.7358874867938e-8
+ k1 = 0.6040969260625 lk1 = -7.0073367568183e-8
+ k2 = 0.019548143337625 lk2 = 1.81509167730435e-8
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 297115.1625125 lvsat = -0.765752570835249
+ ua = 2.45140613429905e-09 lua = 1.99819560766456e-15
+ ub = 2.39982194675e-19 lub = -2.0237801217014e-24 wub = 1.10202595389589e-39 pub = 8.4077907859489e-45
+ uc = -5.150363640875e-11 luc = 9.09268954248117e-17
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.02071299460625 lu0 = 5.24592970319174e-9
+ a0 = 0.912995345534624 la0 = -1.5831450015079e-7
+ keta = -0.004975149172625 lketa = -2.32666555200977e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.1193446512225 lags = 2.06605389098843e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0947667260771126+0*(0.009/sqrt(l*w*mult))} lvoff = 1.2316906862687e-8
+ nfactor = {1.7731568903+0*(0.02/sqrt(l*w*mult))} lnfactor = -5.94283423310471e-8
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.0800000000000101
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.643778489125226 lpclm = 5.73483365645371e-06 wpclm = -1.6940658945086e-21 ppclm = 6.46234853557053e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00454411319014037 lpdiblc2 = -1.26422134731294e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 560706123.996462 lpscbe1 = -1789.84098819564
+ pscbe2 = -1.51292780647975e-08 lpscbe2 = 2.37576760719748e-13 ppscbe2 = 1.54074395550979e-33
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 7.7982685969875e-05 lalpha0 = -2.15382557029979e-10
+ alpha1 = 0.0
+ beta0 = 39.1348639430787 lbeta0 = -6.85062513708628e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 6.543926432625e-09 lagidl = 6.47968046988402e-15
+ bgidl = 1479758789.5 lbgidl = 1773.66032008645
+ cgidl = 931.1572025 lcgidl = -0.00182267338592649
+ egidl = 1.20611845100666 legidl = -4.04192887188653e-6
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.585180250337499 lkt1 = 7.45151766599343e-8
+ kt2 = -0.019032
+ at = 671539.8516375 lat = -1.90454052246243
+ ute = -1.221579087125 lute = -1.29961207391481e-6
+ ua1 = 1.37134480442e-09 lua1 = -5.24182485892768e-15
+ ub1 = -2.61372693375e-18 lub1 = -4.18908547101591e-24
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.11 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 1.5e-05 wmax = 2.0e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.9582756181165+0*(0.0/sqrt(l*w*mult))} lvth0 = -5.65592408254903e-8
+ k1 = 0.6023840567 lk1 = -6.34188786592171e-8
+ k2 = 0.02423914419975 lk2 = -7.35981213077727e-11
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 84741.5405 lvsat = 0.0593178888152024
+ ua = 3.31429591882863e-09 lua = -1.35412689078392e-15
+ ub = -1.22040265805e-18 lub = 3.64980772921096e-24
+ uc = -5.45822372525e-11 luc = 1.02887244309776e-16
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0211909620139 lu0 = 3.38902871430855e-9
+ a0 = 0.823815148711749 la0 = 1.88150118605095e-7
+ keta = -0.00516198539 lketa = -2.25407977497769e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.1427222865525 lags = 1.1578339272997e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0644364973897325+0*(0.009/sqrt(l*w*mult))} lvoff = -1.05515879936641e-7
+ nfactor = {2.19899029989+0*(0.02/sqrt(l*w*mult))} lnfactor = -1.71378900942115e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.01986865950001 leta0 = 2.33609957185798e-7
+ etab = -0.12173557277 letab = 2.00992441533586e-7
+ dsub = 0.811505457875001 ldsub = -9.77097446317086e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.04601663892438 lpclm = -8.30011967043352e-7
+ pdiblc1 = 0.5791285228315 lpdiblc1 = -7.34763365557764e-7
+ pdiblc2 = -0.00110255629368 lpdiblc2 = 9.29506923816533e-9
+ pdiblcb = 0.1634995 lpdiblcb = -7.323196150025e-07 wpdiblcb = -4.2351647362715e-22 ppdiblcb = 3.23117426778526e-27
+ drout = 0.1453011 ldrout = 1.6111031530055e-6
+ pscbe1 = -152915980.78355 lpscbe1 = 982.577320764189 ppscbe1 = 3.46944695195361e-18
+ pscbe2 = 7.56929177375625e-08 lpscbe2 = -1.15267015861442e-13
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 4.37897997750275e-05 lalpha0 = -8.2543365127428e-11
+ alpha1 = -9.424975e-11 lalpha1 = 3.6615980750125e-16
+ beta0 = 69.7665703037275 lbeta0 = -0.000125854651189675
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 9.1846459195e-09 lagidl = -3.7795015330279e-15
+ bgidl = 2611316709.5 lbgidl = -2622.43654132395
+ cgidl = 455.826641375 lcgidl = 2.39834673913322e-5
+ egidl = -1.56307736015895 legidl = 6.71638300851282e-06 wegidl = 6.7762635780344e-21 pegidl = 2.58493941422821e-26
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.5669424975 lkt1 = 3.66159807501186e-9
+ kt2 = -0.019032
+ at = 210065.598725 lat = -0.111715357268631
+ ute = -1.70322385975 lute = 5.71575459509449e-7
+ ua1 = -4.7771419424e-10 lua1 = 1.94176010557143e-15 wua1 = 7.88860905221012e-31 pua1 = 1.50463276905253e-36
+ ub1 = -3.71961517675e-18 lub1 = 1.07284823597862e-25
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.12 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 1.5e-05 wmax = 2.0e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.00534174265973+0*(0.0/sqrt(l*w*mult))} lvth0 = 3.21601686078806e-08 wvth0 = -1.00859244146878e-07 pvth0 = 1.90119170920652e-13
+ k1 = 0.55931480325 lk1 = 1.77664487477661e-8
+ k2 = 0.0190941971058686 lk2 = 9.62460142592328e-09 wk2 = -2.4111688003873e-09 pk2 = 4.54504113288595e-15
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 176673.743395 lvsat = -0.113973853980858
+ ua = 3.43567369390255e-09 lua = -1.58292338990938e-15 wua = -3.8209307616884e-17 pua = 7.20243538113166e-23
+ ub = 1.54521285907453e-18 lub = -1.56336369249119e-24 wub = -1.72100499795403e-23 pub = 3.24408581611836e-29
+ uc = 5.181291727e-13 luc = -9.76670899893637e-19
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.028136701756356 lu0 = -9.70365597152237e-09 wu0 = -3.8884754241122e-08 pu0 = 7.32975673207435e-14
+ a0 = 0.958655606501238 la0 = -6.60234701258035e-08 wa0 = 5.61131674267569e-07 pa0 = -1.05773040033602e-12
+ keta = 0.04266318224 lketa = -1.12690999606489e-07 pketa = 4.03896783473158e-28
+ a1 = 0.0
+ a2 = 0.5
+ ags = -0.34618057285321 lags = 1.03736283819544e-06 wags = 9.07403191879023e-07 pags = -1.710450479676e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.158164876157715+0*(0.009/sqrt(l*w*mult))} lvoff = 7.11616453991121e-08 wvoff = 1.6940658945086e-21
+ nfactor = {1.03301375345643+0*(0.02/sqrt(l*w*mult))} lnfactor = 4.84070950723403e-07 wnfactor = 1.25614975031202e-07 pnfactor = -2.36783599858948e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.4424975e-05 lcit = -8.34105575012501e-12
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.271072766617294 leta0 = -2.39908528709746e-07 weta0 = -7.17389251468121e-10 peta0 = 1.35227515207632e-15
+ etab = -0.02847850446 letab = 2.52033340545777e-8
+ dsub = 0.07100740505 ldsub = 4.18737680767775e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.0769866827459005 lpclm = 9.96604655203293e-7
+ pdiblc1 = 0.00331213796899976 lpdiblc1 = 3.50647640826125e-7
+ pdiblc2 = 0.0058837902087835 lpdiblc2 = -3.87415898724585e-9
+ pdiblcb = -0.401999 lpdiblcb = 3.33642230005e-7
+ drout = 1.52153692559705 ldrout = -9.83094497065812e-07 pdrout = -1.29246970711411e-26
+ pscbe1 = 429292893.4686 lpscbe1 = -114.883496156744
+ pscbe2 = 1.453303481712e-08 lpscbe2 = 1.90576441778914e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -6.0014119919695e-05 lalpha0 = 1.13126504477526e-10 walpha0 = 7.36543649986754e-26 palpha0 = -1.93957696360254e-31
+ alpha1 = 1.884995e-10 lalpha1 = -1.668211150025e-16
+ beta0 = -38.730102860375 lbeta0 = 7.86610352412926e-05 wbeta0 = 1.0842021724855e-19 pbeta0 = -3.6189151799195e-25
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -2.72478415139044e-09 lagidl = 1.86697146034502e-14 wagidl = 1.33258326901749e-13 pagidl = -2.51191279918163e-19
+ bgidl = 1044762109.70235 lbgidl = 330.511046521627 wbgidl = -3598.12386106339 pbgidl = 0.00678244548748513
+ cgidl = 88.0793241694259 lcgidl = 0.000717185321587253 wcgidl = 0.00705147114073484 pcgidl = -1.32919878429295e-8
+ egidl = 3.0805973382958 legidl = -2.03692057970089e-06 wegidl = 2.71050543121376e-20
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.51528141100757 lkt1 = -9.37192916577861e-08 wkt1 = 2.66133421676282e-07 pkt1 = -5.01660169192699e-13
+ kt2 = -0.019032
+ at = 263201.617003028 lat = -0.211876486042623 wat = -0.106453368670515 pat = 2.00664067677075e-7
+ ute = -1.2168945345 lute = -3.45152886940173e-7
+ ua1 = 6.697326371e-10 lua1 = -2.21171434270314e-16
+ ub1 = -3.5355262185e-18 lub1 = -2.39721942258591e-25 wub1 = -4.70197740328915e-38
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.81e-6
+ sbref = 2.81e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.13 pmos
* DC IV MOS Parameters
+ lmin = 8.0e-07 lmax = 1e-06 wmin = 1.5e-05 wmax = 2.0e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.08815164003635+0*(0.0/sqrt(l*w*mult))} lvth0 = 1.05446513736697e-07 wvth0 = 5.04296220734377e-07 pvth0 = -3.45440389721966e-13
+ k1 = 0.589870423500001 lk1 = -9.27512239538251e-9
+ k2 = 0.0147702096506571 lk2 = 1.34513087038482e-08 wk2 = 1.20558440019361e-08 pk2 = -8.2581928621062e-15
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 6575.92405749997 lvsat = 0.0365618656437329
+ ua = -7.46834979143233e-10 lua = 2.11857587319277e-15 wua = 1.91046538084521e-16 pua = -1.30865923355207e-22
+ ub = -2.62100426372647e-19 lub = 3.60995285631332e-26 wub = 8.60502498977017e-23 pub = -5.89439909286762e-29
+ uc = 5.8546574915e-12 luc = -5.69947177939004e-18 wuc = 2.46519032881566e-32 puc = -2.35098870164458e-38
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0106993910442197 lu0 = 5.72827682216467e-09 wu0 = 1.9442377120561e-07 pu0 = -1.33179311156987e-13
+ a0 = 1.0229090794988 la0 = -1.22887472461283e-07 wa0 = -2.8056583713379e-06 pa0 = 1.9218619560746e-12
+ keta = -0.15139736295 lketa = 5.90516125839352e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 1.18515583861605 lags = -3.17862229272805e-07 wags = -4.53701595939514e-06 pags = 3.1078332471059e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0946561577387+0*(0.009/sqrt(l*w*mult))} lvoff = 1.49567471418758e-8
+ nfactor = {0.878622156567864+0*(0.02/sqrt(l*w*mult))} lnfactor = 6.20706742011794e-07 wnfactor = -6.2807487515601e-07 pnfactor = 4.30228149107494e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -1.2124875e-05 lcit = 1.5155428750625e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -0.00024739821325692 leta0 = 2.08460564466848e-10 weta0 = 3.58694625735297e-09 peta0 = -2.4570402515555e-15
+ etab = 0.00072873193075 letab = -6.44924115054096e-10
+ dsub = 1.4666427665 ldsub = -8.16392635938668e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.99390052644125 lpclm = -6.99854511897874e-7
+ pdiblc1 = 0.20282696902275 lpdiblc1 = 1.74078012917712e-7
+ pdiblc2 = -0.0324173066339675 lpdiblc2 = 3.00221202131046e-08 ppdiblc2 = 1.0097419586829e-28
+ pdiblcb = -0.025
+ drout = 0.338402093148499 ldrout = 6.39739139769935e-8
+ pscbe1 = -44797159.5074997 lpscbe1 = 304.68383027684
+ pscbe2 = 1.815406017615e-08 lpscbe2 = -3.18553169343687e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.00024102438742525 lalpha0 = -1.53291069330214e-10
+ alpha1 = 0.0
+ beta0 = 66.614022720125 lbeta0 = -1.4567989176822e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 4.23837552669523e-08 lagidl = -2.1251117239086e-14 wagidl = -6.66291634508747e-13 pagidl = 4.5640643818032e-19
+ bgidl = 85644131.488266 lbgidl = 1179.32566165119 wbgidl = 17990.6193053169 pbgidl = -0.0123234842710455
+ cgidl = 2194.68841540287 lcgidl = -0.00114715319110889 wcgidl = -0.0352573557036742 pcgidl = 2.41511123702384e-8
+ egidl = 1.79942371219525 legidl = -9.03088326470036e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.544732407462151 lkt1 = -6.76553070504645e-08 wkt1 = -1.33066710838144e-06 pkt1 = 9.1150031590573e-13
+ kt2 = -0.019032
+ at = 19653.76998486 lat = 0.00366214082922084 wat = 0.532266843352571 pat = -3.64600126362294e-7
+ ute = -2.0422143225 lute = 3.85250998840887e-7
+ ua1 = -3.42631855000012e-11 lua1 = 4.01861348751573e-16
+ ub1 = -4.5444821125e-18 lub1 = 6.53198979151937e-25
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.41e-6
+ sbref = 2.41e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.14 pmos
* DC IV MOS Parameters
+ lmin = 6e-07 lmax = 8.0e-07 wmin = 1.5e-05 wmax = 2.0e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.881892254404997+0*(0.0/sqrt(l*w*mult))} lvth0 = -3.58401341238471e-8
+ k1 = 0.593523072749999 lk1 = -1.17771688683856e-8
+ k2 = 0.0189560867924999 lk2 = 1.05840037910714e-8
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 61502.5565075001 lvsat = -0.00106260295135502
+ ua = -1.82337677780051e-09 lua = 2.85600162256401e-15
+ ub = 2.469434477865e-18 lub = -1.83498822316514e-24 wub = 1.17549435082229e-38 pub = -8.4077907859489e-45
+ uc = 2.53255847000001e-12 luc = -3.42385056015765e-18
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.00709052591749998 lu0 = 8.20033138964208e-9
+ a0 = 0.93451931175 la0 = -6.2340923502192e-8
+ keta = 0.0117180821250003 lketa = -5.26816517152144e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = -0.561400778000003 lags = 8.7852032032611e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {0.00731538466477499+0*(0.009/sqrt(l*w*mult))} lvoff = -5.48932495467926e-8
+ nfactor = {1.78668573025+0*(0.02/sqrt(l*w*mult))} lnfactor = -1.31226564259923e-9
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -0.0573036120981399 leta0 = 3.92916817945423e-08 weta0 = 1.7205356741103e-22 peta0 = -1.89326617253043e-29
+ etab = -0.00072873193075 letab = 3.53431342754096e-10
+ dsub = 0.193392103971499 ldsub = 5.57777016400423e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.25744420752125 lpclm = 4.89609384280731e-7
+ pdiblc1 = 0.189717426328749 lpdiblc1 = 1.83057984115388e-7
+ pdiblc2 = 0.02598707339889 lpdiblc2 = -9.98458808750265e-9
+ pdiblcb = -0.025
+ drout = -0.682593035841502 ldrout = 7.63350472359499e-7
+ pscbe1 = 430689610.608999 lpscbe1 = -21.0222298191115
+ pscbe2 = 1.0686514267575e-08 lpscbe2 = 1.92969991620746e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -0.000115023676316125 lalpha0 = 9.06000740923091e-11 palpha0 = 1.97215226305253e-31
+ alpha1 = 0.0
+ beta0 = 27.36521542835 lbeta0 = 1.23172475740074e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 2.30942115275e-08 lagidl = -8.03787622527987e-15
+ bgidl = 2050039997.49999 lbgidl = -166.275684587514
+ cgidl = 1223.24275 lcgidl = -0.00048171776753625
+ egidl = -0.212081994370002 legidl = 4.74783024998628e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.704172874499999 lkt1 = 4.15606156681274e-8
+ kt2 = -0.019032
+ at = 41974.825 lat = -0.011627670250875
+ ute = -1.6071111875 lute = 8.72075268815616e-8
+ ua1 = 5.53369989999999e-10 lua1 = -6.64438300049995e-19
+ ub1 = -4.2982652075e-18 lub1 = 4.8454163031146e-25
+ uc1 = -2.733805074e-10 luc1 = 1.12462826666463e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.02e-6
+ sbref = 2.01e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.15 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 6e-07 wmin = 1.5e-05 wmax = 2.0e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.724081721364389+0*(0.0/sqrt(l*w*mult))} lvth0 = -1.12377453595879e-07 wvth0 = -2.78060744401552e-06 pvth0 = 1.3485807073103e-12
+ k1 = 0.458361439999999 lk1 = 5.37755472071992e-8
+ k2 = 0.0598778056171021 lk2 = -9.26282523026648e-09 wk2 = -3.83908927875429e-07 pk2 = 1.86193910474944e-13
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 48942.9706761565 lvsat = 0.00502873337891746 wvsat = -0.204272892745298 pvsat = 9.90713316170058e-8
+ ua = 1.1403463188889e-08 lua = -3.55894962708056e-15 wua = 7.74046534978503e-17 pua = -3.754086992322e-23
+ ub = -6.50578006718928e-18 lub = 2.51794595511346e-24 wub = -1.89754744507789e-23 pub = 9.20301023125551e-30
+ uc = -1.622212725e-12 luc = -1.40880730443863e-18
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0401817739318384 lu0 = -7.84875844107197e-09 wu0 = -4.95284195853768e-08 pu0 = 2.40210358568097e-14
+ a0 = 0.214396682999999 la0 = 2.86914950828416e-7
+ keta = -0.13938919825 lketa = 2.06046237302588e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 1.25
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1225417579515+0*(0.009/sqrt(l*w*mult))} lvoff = 8.08681533638781e-9
+ nfactor = {-1.93227371694453+0*(0.02/sqrt(l*w*mult))} lnfactor = 1.80236447144951e-06 wnfactor = 6.46092328981187e-05 pnfactor = -3.13351549094231e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 2.924975e-05 lcit = -9.33603250125001e-12
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -0.32283809676168 leta0 = 1.68074579183936e-07 weta0 = 2.59520582848481e-06 peta0 = -1.25866185078599e-12
+ etab = 0.014823462485 letab = -7.18930518791258e-9
+ dsub = 0.419003534557 ldsub = -5.36427141367725e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.998842207074997 lpclm = 1.3003506148716e-7
+ pdiblc1 = 1.618697765494 lpdiblc1 = -5.09990335478063e-7
+ pdiblc2 = 0.00770696779004999 lpdiblc2 = -1.1188282677433e-9
+ pdiblcb = -0.025
+ drout = 0.859530092143 ldrout = 1.5428465902656e-8
+ pscbe1 = 482455064.779999 lpscbe1 = -46.1282162647763
+ pscbe2 = 1.53528728706e-08 lpscbe2 = -3.33460674466638e-16
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -2.58245787588002e-05 lalpha0 = 4.73389577724941e-11
+ alpha1 = 0.0
+ beta0 = 45.3597691823499 lbeta0 = 3.5899789760862e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -2.43855339383308e-08 lagidl = 1.49895629269208e-14 wagidl = 5.09408710088021e-14 pagidl = -2.47060677349141e-20
+ bgidl = 2121918485.0757 lbgidl = -201.13639166929 wbgidl = -1157.74706838187 pbgidl = 0.000561501539429854
+ cgidl = -8725.95252414812 lcgidl = 0.00434359219444922 wcgidl = 0.12951021805747 pcgidl = -6.28118082067826e-8
+ egidl = 1.15799168033 legidl = -1.89695856862498e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.5220735098486 lkt1 = -4.67566656909789e-08 wkt1 = -2.31549413676373e-06 pkt1 = 1.12300307885973e-12
+ kt2 = -0.019032
+ at = 18000.0
+ ute = -1.638662255 lute = 1.02509636863726e-7
+ ua1 = 5.52e-10
+ ub1 = -7.68506303999999e-18 lub1 = 2.1271216450848e-24
+ uc1 = -4.1496e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 1.81e-6
+ sbref = 1.81e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.16 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 1.0e-05 wmax = 1.5e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.979018+0*(0.0/sqrt(l*w*mult))}
+ k1 = 0.59521
+ k2 = 0.0218501
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200000.0
+ ua = 2.70482362e-9
+ ub = -1.668e-20
+ uc = -3.9972e-11
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0213783
+ a0 = 0.8929174
+ keta = -0.0079259
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.145547
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.093204657+0*(0.009/sqrt(l*w*mult))}
+ nfactor = {1.76562+0*(0.02/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.0800000000000101
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.08353125
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0029407877
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 333712830.0
+ pscbe2 = 1.5000958e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 5.0667189e-5
+ alpha1 = 0.0
+ beta0 = 38.266046
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 7.3657e-9
+ bgidl = 1704700000.0
+ cgidl = 700.0
+ egidl = 0.69350825
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.57573
+ kt2 = -0.019032
+ at = 430000.0
+ ute = -1.3864
+ ua1 = 7.0656e-10
+ ub1 = -3.145e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.17 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 1.0e-05 wmax = 1.5e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.979018+0*(0.0/sqrt(l*w*mult))}
+ k1 = 0.59521
+ k2 = 0.0218501
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200000.0
+ ua = 2.70482362e-9
+ ub = -1.668e-20
+ uc = -3.9972e-11
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0213783
+ a0 = 0.8929174
+ keta = -0.0079259
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.145547
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.093204657+0*(0.009/sqrt(l*w*mult))}
+ nfactor = {1.76562+0*(0.02/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.0800000000000101
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.08353125
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0029407877
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 333712830.0
+ pscbe2 = 1.5000958e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 5.0667189e-5
+ alpha1 = 0.0
+ beta0 = 38.266046
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 7.3657e-9
+ bgidl = 1704700000.0
+ cgidl = 700.0
+ egidl = 0.69350825
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.57573
+ kt2 = -0.019032
+ at = 430000.0
+ ute = -1.3864
+ ua1 = 7.0656e-10
+ ub1 = -3.145e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.18 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 1.0e-05 wmax = 1.5e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.985024202270001+0*(0.0/sqrt(l*w*mult))} lvth0 = 4.73588748679414e-8
+ k1 = 0.6040969260625 lk1 = -7.0073367568183e-8
+ k2 = 0.019548143337625 lk2 = 1.81509167730436e-8
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 297115.1625125 lvsat = -0.76575257083525 wvsat = 1.77635683940025e-15
+ ua = 2.45140613429905e-09 lua = 1.99819560766456e-15
+ ub = 2.39982194675e-19 lub = -2.0237801217014e-24 wub = -3.67341984631965e-40 pub = -2.10194769648723e-45
+ uc = -5.150363640875e-11 luc = 9.09268954248117e-17
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.02071299460625 lu0 = 5.24592970319185e-9
+ a0 = 0.912995345534624 la0 = -1.5831450015079e-7
+ keta = -0.004975149172625 lketa = -2.32666555200977e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.1193446512225 lags = 2.06605389098844e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0947667260771126+0*(0.009/sqrt(l*w*mult))} lvoff = 1.23169068626865e-8
+ nfactor = {1.7731568903+0*(0.02/sqrt(l*w*mult))} lnfactor = -5.94283423310471e-8
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.0800000000000101
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.643778489125225 lpclm = 5.7348336564537e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00454411319014037 lpdiblc2 = -1.26422134731294e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 560706123.996463 lpscbe1 = -1789.84098819564 wpscbe1 = -3.63797880709171e-12
+ pscbe2 = -1.51292780647975e-08 lpscbe2 = 2.37576760719748e-13 ppscbe2 = 3.85185988877447e-34
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 7.7982685969875e-05 lalpha0 = -2.1538255702998e-10
+ alpha1 = 0.0
+ beta0 = 39.1348639430787 lbeta0 = -6.85062513708628e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 6.543926432625e-09 lagidl = 6.47968046988405e-15
+ bgidl = 1479758789.5 lbgidl = 1773.66032008645
+ cgidl = 931.1572025 lcgidl = -0.00182267338592649
+ egidl = 1.20611845100666 legidl = -4.04192887188653e-6
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.5851802503375 lkt1 = 7.45151766599359e-8
+ kt2 = -0.019032
+ at = 671539.8516375 lat = -1.90454052246243
+ ute = -1.221579087125 lute = -1.29961207391482e-6
+ ua1 = 1.37134480442e-09 lua1 = -5.24182485892768e-15
+ ub1 = -2.61372693375e-18 lub1 = -4.18908547101592e-24
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.19 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 1.0e-05 wmax = 1.5e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.9582756181165+0*(0.0/sqrt(l*w*mult))} lvth0 = -5.65592408254869e-8
+ k1 = 0.6023840567 lk1 = -6.34188786592163e-8
+ k2 = 0.02423914419975 lk2 = -7.35981213077727e-11
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 84741.5405 lvsat = 0.0593178888152022
+ ua = 3.31429591882862e-09 lua = -1.35412689078391e-15
+ ub = -1.22040265805e-18 lub = 3.64980772921096e-24 wub = 2.93873587705572e-39
+ uc = -5.45822372525e-11 luc = 1.02887244309776e-16
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0211909620139 lu0 = 3.38902871430855e-9
+ a0 = 0.82381514871175 la0 = 1.88150118605095e-7
+ keta = -0.00516198539000001 lketa = -2.2540797749777e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.1427222865525 lags = 1.1578339272997e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0644364973897326+0*(0.009/sqrt(l*w*mult))} lvoff = -1.05515879936641e-7
+ nfactor = {2.19899029989+0*(0.02/sqrt(l*w*mult))} lnfactor = -1.71378900942115e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.0198686595000101 leta0 = 2.33609957185798e-7
+ etab = -0.12173557277 letab = 2.00992441533586e-7
+ dsub = 0.811505457875 ldsub = -9.77097446317087e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.04601663892437 lpclm = -8.30011967043354e-7
+ pdiblc1 = 0.5791285228315 lpdiblc1 = -7.34763365557764e-07 wpdiblc1 = -3.3881317890172e-21
+ pdiblc2 = -0.00110255629368 lpdiblc2 = 9.29506923816533e-9
+ pdiblcb = 0.1634995 lpdiblcb = -7.323196150025e-07 ppdiblcb = 8.07793566946316e-28
+ drout = 0.1453011 ldrout = 1.6111031530055e-6
+ pscbe1 = -152915980.78355 lpscbe1 = 982.577320764188
+ pscbe2 = 7.56929177375625e-08 lpscbe2 = -1.15267015861442e-13
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 4.37897997750275e-05 lalpha0 = -8.2543365127428e-11
+ alpha1 = -9.424975e-11 lalpha1 = 3.6615980750125e-16
+ beta0 = 69.7665703037275 lbeta0 = -0.000125854651189675
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 9.1846459195e-09 lagidl = -3.7795015330279e-15
+ bgidl = 2611316709.5 lbgidl = -2622.43654132395 wbgidl = 1.45519152283669e-11
+ cgidl = 455.826641375 lcgidl = 2.39834673913322e-5
+ egidl = -1.56307736015895 legidl = 6.71638300851282e-06 pegidl = 3.23117426778526e-27
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.5669424975 lkt1 = 3.6615980750127e-9
+ kt2 = -0.019032
+ at = 210065.598725 lat = -0.111715357268631
+ ute = -1.70322385975 lute = 5.71575459509449e-7
+ ua1 = -4.7771419424e-10 lua1 = 1.94176010557143e-15 wua1 = 5.91645678915759e-31 pua1 = -1.1284745767894e-36
+ ub1 = -3.71961517675e-18 lub1 = 1.07284823597868e-25
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.20 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 1.0e-05 wmax = 1.5e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.979524856972231+0*(0.0/sqrt(l*w*mult))} lvth0 = -1.65045318286305e-08 wvth0 = -4.88641414179582e-07 pvth0 = 9.21086622521448e-13
+ k1 = 0.55931480325 lk1 = 1.77664487477661e-8
+ k2 = 0.0188714178323469 lk2 = 1.00445392426153e-08 wk2 = 9.35084158635998e-10 pk2 = -1.76262896360825e-15
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 176673.743395 lvsat = -0.113973853980858
+ ua = 3.43253664181811e-09 lua = -1.57701006241549e-15 wua = 8.91073929857826e-18 pua = -1.67966990241309e-23
+ ub = -2.5387930966269e-19 lub = 1.82791605011762e-24 wub = 9.8131887536867e-24 pub = -1.84978117347557e-29
+ uc = 5.181291727e-13 luc = -9.76670899893637e-19
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0221875388346815 lu0 = 1.51048639001957e-09 wu0 = 5.04745641356098e-08 pu0 = -9.51443010228038e-14
+ a0 = 0.992705570208177 la0 = -1.3020748146356e-07 wa0 = 4.96846711070198e-08 pa0 = -9.36553566133752e-14
+ keta = 0.04266318224 lketa = -1.12690999606489e-07 pketa = 2.01948391736579e-28
+ a1 = 0.0
+ a2 = 0.5
+ ags = -0.291044266088503 lags = 9.33431175625497e-07 wags = 7.92290680280283e-08 pags = -1.49346397087494e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.158164876157715+0*(0.009/sqrt(l*w*mult))} lvoff = 7.1161645399112e-8
+ nfactor = {1.32338160786073+0*(0.02/sqrt(l*w*mult))} lnfactor = -6.32710029894297e-08 wnfactor = -4.23585131689861e-06 pnfactor = 7.98455855309729e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.4424975e-05 lcit = -8.34105575012501e-12
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.271025005895605 leta0 = -2.39818499988167e-7
+ etab = -0.02847850446 letab = 2.52033340545777e-8
+ dsub = 0.07100740505 ldsub = 4.18737680767775e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.077008852945919 lpclm = 9.96562864487108e-07 wpclm = -3.33007179001573e-10 ppclm = 6.27716867386064e-16
+ pdiblc1 = 0.00331213796899998 lpdiblc1 = 3.50647640826125e-7
+ pdiblc2 = 0.0058837902087835 lpdiblc2 = -3.87415898724585e-09 wpdiblc2 = -2.64697796016969e-23
+ pdiblcb = -0.401999 lpdiblcb = 3.33642230005e-7
+ drout = 1.52153692559705 ldrout = -9.83094497065811e-7
+ pscbe1 = 429292893.4686 lpscbe1 = -114.883496156744
+ pscbe2 = 1.453303481712e-08 lpscbe2 = 1.90576441778787e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -6.0014119919695e-05 lalpha0 = 1.13126504477525e-10 walpha0 = 7.67814096269715e-26 palpha0 = 1.42007993059562e-31
+ alpha1 = 1.884995e-10 lalpha1 = -1.668211150025e-16
+ beta0 = -38.730102860375 lbeta0 = 7.86610352412926e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 6.146987834e-09 lagidl = 1.94646876984916e-15
+ bgidl = 805214344.0 lbgidl = 782.05738713172
+ cgidl = 557.53624725 lcgidl = -0.000167738631135014 wcgidl = -3.46944695195361e-18
+ egidl = 3.0805973382958 legidl = -2.03692057970089e-06 wegidl = 1.35525271560688e-20 pegidl = 1.29246970711411e-26
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.477698881783043 lkt1 = -1.64562171333373e-07 wkt1 = -2.98374432385308e-07 pkt1 = 5.62434313174146e-13
+ kt2 = -0.019032
+ at = 252921.896197275 lat = -0.192499263722382 wat = 0.04795303377621 pat = -9.03912289029879e-8
+ ute = -0.957769236678804 lute = -8.33602777706637e-07 wute = -3.8921879081691e-06 pute = 7.3367547459592e-12
+ ua1 = 9.04878646580727e-10 lua1 = -6.64420486411436e-16 wua1 = -3.53200734336112e-15 pua1 = 6.65781618219899e-21
+ ub1 = -3.15331197017373e-18 lub1 = -9.60193889282366e-25 wub1 = -5.74104376598523e-24 pub1 = 1.08218387936633e-29
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.81e-6
+ sbref = 2.81e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.21 pmos
* DC IV MOS Parameters
+ lmin = 8.0e-07 lmax = 1e-06 wmin = 1.0e-05 wmax = 1.5e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.21723606847385+0*(0.0/sqrt(l*w*mult))} lvth0 = 1.93868701794243e-07 wvth0 = 2.44320707089792e-06 pvth0 = -1.67358462752972e-12
+ k1 = 0.5898704235 lk1 = -9.27512239538167e-9
+ k2 = 0.0158841060182657 lk2 = 1.2688295261518e-08 wk2 = -4.67542079318063e-09 pk2 = 3.20263986622459e-15
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 6575.92405749997 lvsat = 0.0365618656437328
+ ua = -7.31149718721071e-10 lua = 2.10783154822989e-15 wua = -4.45536964929418e-17 pua = 3.05190593291869e-23
+ ub = 8.73336041731344e-18 lub = -6.12574617205763e-24 wub = -4.90659437684335e-23 pub = 3.36099261516581e-29
+ uc = 5.8546574915e-12 luc = -5.69947177939004e-18 wuc = -1.23259516440783e-32
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0404452056525925 lu0 = -1.46474574554976e-08 wu0 = -2.52372820678049e-07 pu0 = 1.7287412030036e-13
+ a0 = 0.852659260964119 la0 = -6.26719801411757e-09 wa0 = -2.48423355535092e-07 pa0 = 1.70168756424763e-13
+ keta = -0.15139736295 lketa = 5.90516125839353e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.909474304792512 lags = -1.29021757011348e-07 wags = -3.96145340140152e-07 pags = 2.71357577269294e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0946561577386997+0*(0.009/sqrt(l*w*mult))} lvoff = 1.49567471418758e-8
+ nfactor = {-0.57321711545363+0*(0.02/sqrt(l*w*mult))} lnfactor = 1.61520938415016e-06 wnfactor = 2.1179256584493e-05 pnfactor = -1.45076848640948e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -1.2124875e-05 lcit = 1.5155428750625e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -8.59460481489999e-06 leta0 = 4.48812867021009e-11
+ etab = 0.00072873193075 letab = -6.44924115054096e-10
+ dsub = 1.4666427665 ldsub = -8.16392635938667e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.99378967544115 lpclm = -6.99778579517064e-07 wpclm = 1.66503589502142e-09 ppclm = -1.14054126290564e-15
+ pdiblc1 = 0.20282696902275 lpdiblc1 = 1.74078012917712e-7
+ pdiblc2 = -0.0324173066339675 lpdiblc2 = 3.00221202131046e-08 wpdiblc2 = -7.94093388050907e-23 ppdiblc2 = 2.52435489670724e-29
+ pdiblcb = -0.025
+ drout = 0.338402093148499 ldrout = 6.39739139769931e-8
+ pscbe1 = -44797159.5074997 lpscbe1 = 304.68383027684
+ pscbe2 = 1.815406017615e-08 lpscbe2 = -3.18553169343687e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.00024102438742525 lalpha0 = -1.53291069330214e-10
+ alpha1 = 0.0
+ beta0 = 66.6140227201249 lbeta0 = -1.4567989176822e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -1.97510466e-09 lagidl = 9.1344800165767e-15
+ bgidl = 1283382960 lbgidl = 358.880552814799
+ cgidl = -152.5962 lcgidl = 0.000460725034019
+ egidl = 1.79942371219525 legidl = -9.03088326470036e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.732645053584783 lkt1 = 6.106391598031e-08 wkt1 = 1.49187216192654e-06 pkt1 = -1.02192497155888e-12
+ kt2 = -0.019032
+ at = 71052.374013626 lat = -0.0315456459374638 wat = -0.239765168881053 pat = 1.64237941857677e-7
+ ute = -3.33784081160598 lute = 1.27274866574604e-06 wute = 1.94609395408455e-05 pute = -1.33306462807814e-11
+ ua1 = -1.20999323290363e-09 lua1 = 1.20723055257282e-15 wua1 = 1.76600367168056e-14 pua1 = -1.20970368508282e-20
+ ub1 = -6.45555335413133e-18 lub1 = 1.96227322431319e-24 wub1 = 2.87052188299261e-23 pub1 = -1.96629313724053e-29
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.41e-6
+ sbref = 2.41e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.22 pmos
* DC IV MOS Parameters
+ lmin = 6e-07 lmax = 8.0e-07 wmin = 1.0e-05 wmax = 1.5e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.881892254405001+0*(0.0/sqrt(l*w*mult))} lvth0 = -3.58401341238471e-8
+ k1 = 0.59352307275 lk1 = -1.1777168868386e-8
+ k2 = 0.0189560867925 lk2 = 1.05840037910715e-8
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 61502.5565075 lvsat = -0.00106260295135502
+ ua = -1.8233767778005e-09 lua = 2.85600162256401e-15
+ ub = 2.469434477865e-18 lub = -1.83498822316514e-24 wub = -2.93873587705572e-39
+ uc = 2.53255847e-12 luc = -3.42385056015765e-18
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.00709052591749998 lu0 = 8.20033138964208e-9
+ a0 = 0.93451931175 la0 = -6.23409235021911e-8
+ keta = 0.011718082125 lketa = -5.26816517152144e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = -0.561400777999999 lags = 8.78520320326111e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {0.00731538466477488+0*(0.009/sqrt(l*w*mult))} lvoff = -5.48932495467926e-8
+ nfactor = {1.78668573025+0*(0.02/sqrt(l*w*mult))} lnfactor = -1.31226564259754e-9
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -0.0573036120981399 leta0 = 3.92916817945423e-08 weta0 = 8.27180612553028e-23 peta0 = 6.7053176943786e-30
+ etab = -0.00072873193075 letab = 3.53431342754096e-10
+ dsub = 0.1933921039715 ldsub = 5.57777016400425e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.257444207521248 lpclm = 4.89609384280732e-7
+ pdiblc1 = 0.18971742632875 lpdiblc1 = 1.83057984115388e-7
+ pdiblc2 = 0.02598707339889 lpdiblc2 = -9.98458808750266e-9
+ pdiblcb = -0.025
+ drout = -0.6825930358415 ldrout = 7.63350472359499e-7
+ pscbe1 = 430689610.609 lpscbe1 = -21.0222298191118
+ pscbe2 = 1.0686514267575e-08 lpscbe2 = 1.92969991620747e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -0.000115023676316125 lalpha0 = 9.06000740923091e-11 palpha0 = 9.86076131526265e-32
+ alpha1 = 0.0
+ beta0 = 27.36521542835 lbeta0 = 1.23172475740074e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 2.30942115275e-08 lagidl = -8.03787622527987e-15
+ bgidl = 2050039997.5 lbgidl = -166.27568458751
+ cgidl = 1223.24275 lcgidl = -0.00048171776753625 wcgidl = 6.93889390390723e-18
+ egidl = -0.212081994370001 legidl = 4.74783024998628e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.704172874499999 lkt1 = 4.15606156681274e-8
+ kt2 = -0.019032
+ at = 41974.825 lat = -0.011627670250875
+ ute = -1.6071111875 lute = 8.72075268815624e-8
+ ua1 = 5.5336999e-10 lua1 = -6.644383000496e-19
+ ub1 = -4.2982652075e-18 lub1 = 4.8454163031146e-25
+ uc1 = -2.733805074e-10 luc1 = 1.12462826666463e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.02e-6
+ sbref = 2.01e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.23 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 6e-07 wmin = 1.0e-05 wmax = 1.5e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.919611169286423+0*(0.0/sqrt(l*w*mult))} lvth0 = -1.75466490009304e-08 wvth0 = 1.56339891085183e-07 pvth0 = -7.58240654768654e-14
+ k1 = 0.45836144 lk1 = 5.37755472072005e-8
+ k2 = 0.0272435108281166 lk2 = 6.56464457091756e-09 wk2 = 1.062740401224e-07 pk2 = -5.15423780891639e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 39223.5637422139 lvsat = 0.00974259714484493 wvsat = -0.0582826769657103 pvsat = 2.82668069149848e-8
+ ua = 1.14039924576892e-08 lua = -3.55920631980234e-15 wua = 6.94547788934178e-17 pua = -3.36852204894646e-23
+ ub = -9.66012090210066e-18 lub = 4.04778548834131e-24 wub = 2.84042578992359e-23 pub = -1.37759230598399e-29
+ uc = -1.622212725e-12 luc = -1.40880730443863e-18
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0309795773262133 lu0 = -3.38573909832685e-09 wu0 = 8.86930456986626e-08 pu0 = -4.30156836986229e-14
+ a0 = 0.214396682999999 la0 = 2.86914950828415e-7
+ keta = -0.13938919825 lketa = 2.06046237302589e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 1.25
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1225417579515+0*(0.009/sqrt(l*w*mult))} lvoff = 8.0868153363877e-9
+ nfactor = {5.13389137034511+0*(0.02/sqrt(l*w*mult))} lnfactor = -1.62469026506053e-06 wnfactor = -4.1528000869204e-05 pnfactor = 2.01408727815596e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 2.924975e-05 lcit = -9.33603250125e-12
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -0.187118725494707 leta0 = 1.02251362716311e-07 weta0 = 5.56634912440451e-07 peta0 = -2.69965149359056e-13
+ etab = -0.0119136626796646 letab = 5.77806683132394e-09 wetab = 4.01604614216093e-07 petab = -1.94776229871734e-13
+ dsub = 0.419003534557 ldsub = -5.36427141367723e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.174036654856533 lpclm = 5.30061630285354e-07 wpclm = 1.23889802498197e-05 ppclm = -6.00859347626132e-12
+ pdiblc1 = 1.618697765494 lpdiblc1 = -5.09990335478062e-7
+ pdiblc2 = 0.00770696779005001 lpdiblc2 = -1.11882826774331e-9
+ pdiblcb = -0.025
+ drout = 0.859530092143002 ldrout = 1.5428465902656e-8
+ pscbe1 = 482455064.78 lpscbe1 = -46.1282162647763
+ pscbe2 = 1.53528728706e-08 lpscbe2 = -3.33460674466651e-16
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -2.58245787588e-05 lalpha0 = 4.73389577724943e-11
+ alpha1 = 0.0
+ beta0 = 45.35976918235 lbeta0 = 3.58997897608609e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -6.85843849803835e-08 lagidl = 3.64257846880611e-14 wagidl = 7.1482909430204e-13 pagidl = -3.46688536591018e-19
+ bgidl = 1564154123.85678 lbgidl = 69.3765347000808 wbgidl = 7220.14471060588 pbgidl = -0.00350173408392031
+ cgidl = -506.471849590308 lcgidl = 0.000357185164692051 wcgidl = 0.00604962365800364 pcgidl = -2.93403722601348e-9
+ egidl = 1.15799168033 legidl = -1.89695856862498e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.676229249999999 lkt1 = 2.800809750375e-8
+ kt2 = -0.019032
+ at = 18000.0
+ ute = -1.638662255 lute = 1.02509636863725e-7
+ ua1 = 5.52e-10
+ ub1 = -7.68506304000001e-18 lub1 = 2.1271216450848e-24
+ uc1 = -4.1496e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 1.81e-6
+ sbref = 1.81e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.24 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 7e-06 wmax = 1.0e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.979018+0*(0.0/sqrt(l*w*mult))}
+ k1 = 0.59521
+ k2 = 0.0218501
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200000.0
+ ua = 2.70482362e-9
+ ub = -1.668e-20
+ uc = -3.9972e-11
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0213783
+ a0 = 0.8929174
+ keta = -0.0079259
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.145547
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.093204657+0*(0.009/sqrt(l*w*mult))}
+ nfactor = {1.76562+0*(0.02/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.0800000000000101
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.08353125
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0029407877
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 333712830.0
+ pscbe2 = 1.5000958e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 5.0667189e-5
+ alpha1 = 0.0
+ beta0 = 38.266046
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 7.3657e-9
+ bgidl = 1704700000.0
+ cgidl = 700.0
+ egidl = 0.69350825
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.57573
+ kt2 = -0.019032
+ at = 430000.0
+ ute = -1.3864
+ ua1 = 7.0656e-10
+ ub1 = -3.145e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.25 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 7e-06 wmax = 1.0e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.979018+0*(0.0/sqrt(l*w*mult))}
+ k1 = 0.59521
+ k2 = 0.0218501
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200000.0
+ ua = 2.70482362e-9
+ ub = -1.668e-20
+ uc = -3.9972e-11
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0213783
+ a0 = 0.8929174
+ keta = -0.0079259
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.145547
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.093204657+0*(0.009/sqrt(l*w*mult))}
+ nfactor = {1.76562+0*(0.02/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.0800000000000101
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.08353125
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0029407877
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 333712830.0
+ pscbe2 = 1.5000958e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 5.0667189e-5
+ alpha1 = 0.0
+ beta0 = 38.266046
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 7.3657e-9
+ bgidl = 1704700000.0
+ cgidl = 700.0
+ egidl = 0.69350825
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.57573
+ kt2 = -0.019032
+ at = 430000.0
+ ute = -1.3864
+ ua1 = 7.0656e-10
+ ub1 = -3.145e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.26 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 7e-06 wmax = 1.0e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.985024202270001+0*(0.0/sqrt(l*w*mult))} lvth0 = 4.73588748679346e-8
+ k1 = 0.6040969260625 lk1 = -7.0073367568183e-8
+ k2 = 0.019548143337625 lk2 = 1.81509167730436e-8
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 297115.1625125 lvsat = -0.76575257083525
+ ua = 2.45140613429905e-09 lua = 1.99819560766457e-15
+ ub = 2.39982194675e-19 lub = -2.0237801217014e-24 wub = -9.18354961579912e-41 pub = -1.75162308040602e-45
+ uc = -5.150363640875e-11 luc = 9.09268954248117e-17
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.02071299460625 lu0 = 5.24592970319185e-9
+ a0 = 0.912995345534625 la0 = -1.5831450015079e-7
+ keta = -0.00497514917262501 lketa = -2.32666555200977e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.1193446512225 lags = 2.06605389098843e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0947667260771126+0*(0.009/sqrt(l*w*mult))} lvoff = 1.2316906862687e-8
+ nfactor = {1.7731568903+0*(0.02/sqrt(l*w*mult))} lnfactor = -5.94283423310538e-8
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.0800000000000101
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.643778489125225 lpclm = 5.7348336564537e-06 wpclm = -8.470329472543e-22
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00454411319014037 lpdiblc2 = -1.26422134731294e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 560706123.996463 lpscbe1 = -1789.84098819564
+ pscbe2 = -1.51292780647975e-08 lpscbe2 = 2.37576760719748e-13
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 7.7982685969875e-05 lalpha0 = -2.1538255702998e-10
+ alpha1 = 0.0
+ beta0 = 39.1348639430788 lbeta0 = -6.85062513708628e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 6.54392643262501e-09 lagidl = 6.47968046988405e-15
+ bgidl = 1479758789.5 lbgidl = 1773.66032008646
+ cgidl = 931.1572025 lcgidl = -0.00182267338592649
+ egidl = 1.20611845100666 legidl = -4.04192887188653e-6
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.5851802503375 lkt1 = 7.45151766599343e-8
+ kt2 = -0.019032
+ at = 671539.8516375 lat = -1.90454052246243
+ ute = -1.221579087125 lute = -1.29961207391481e-6
+ ua1 = 1.37134480442e-09 lua1 = -5.24182485892768e-15
+ ub1 = -2.61372693375e-18 lub1 = -4.18908547101592e-24
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.27 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 7e-06 wmax = 1.0e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.958275618116502+0*(0.0/sqrt(l*w*mult))} lvth0 = -5.65592408254886e-8
+ k1 = 0.602384056700001 lk1 = -6.34188786592171e-8
+ k2 = 0.02423914419975 lk2 = -7.35981213077727e-11
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 84741.5405 lvsat = 0.0593178888152024
+ ua = 3.31429591882862e-09 lua = -1.35412689078392e-15
+ ub = -1.22040265805e-18 lub = 3.64980772921096e-24 wub = 1.46936793852786e-39
+ uc = -5.45822372525e-11 luc = 1.02887244309776e-16
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0211909620139 lu0 = 3.3890287143086e-9
+ a0 = 0.82381514871175 la0 = 1.88150118605095e-7
+ keta = -0.00516198539 lketa = -2.2540797749777e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.1427222865525 lags = 1.15783392729971e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0644364973897326+0*(0.009/sqrt(l*w*mult))} lvoff = -1.05515879936641e-7
+ nfactor = {2.19899029989+0*(0.02/sqrt(l*w*mult))} lnfactor = -1.71378900942115e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.0198686595000102 leta0 = 2.33609957185797e-7
+ etab = -0.12173557277 letab = 2.00992441533586e-7
+ dsub = 0.811505457875 ldsub = -9.77097446317087e-07 wdsub = 3.3881317890172e-21
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.04601663892438 lpclm = -8.30011967043352e-7
+ pdiblc1 = 0.5791285228315 lpdiblc1 = -7.34763365557764e-7
+ pdiblc2 = -0.00110255629368 lpdiblc2 = 9.29506923816534e-09 ppdiblc2 = 1.26217744835362e-29
+ pdiblcb = 0.1634995 lpdiblcb = -7.323196150025e-07 wpdiblcb = 4.2351647362715e-22 ppdiblcb = 4.03896783473158e-28
+ drout = 0.1453011 ldrout = 1.6111031530055e-6
+ pscbe1 = -152915980.78355 lpscbe1 = 982.577320764188 ppscbe1 = -1.73472347597681e-18
+ pscbe2 = 7.56929177375625e-08 lpscbe2 = -1.15267015861442e-13
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 4.37897997750275e-05 lalpha0 = -8.2543365127428e-11
+ alpha1 = -9.42497499999999e-11 lalpha1 = 3.6615980750125e-16
+ beta0 = 69.7665703037275 lbeta0 = -0.000125854651189675
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 9.1846459195e-09 lagidl = -3.7795015330279e-15
+ bgidl = 2611316709.5 lbgidl = -2622.43654132395
+ cgidl = 455.826641375 lcgidl = 2.39834673913314e-5
+ egidl = -1.56307736015895 legidl = 6.71638300851282e-06 pegidl = -8.07793566946316e-27
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.5669424975 lkt1 = 3.66159807501186e-9
+ kt2 = -0.019032
+ at = 210065.598725 lat = -0.111715357268632
+ ute = -1.70322385975 lute = 5.71575459509453e-7
+ ua1 = -4.7771419424e-10 lua1 = 1.94176010557143e-15 wua1 = -7.88860905221012e-31 pua1 = -7.52316384526264e-37
+ ub1 = -3.71961517675e-18 lub1 = 1.07284823597868e-25
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.28 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 7e-06 wmax = 1.0e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.028289099962+0*(0.0/sqrt(l*w*mult))} lvth0 = 7.54158223858703e-8
+ k1 = 0.55931480325 lk1 = 1.77664487477661e-8
+ k2 = 0.0189647350785 lk2 = 9.86863670020288e-9
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 176673.743395 lvsat = -0.113973853980858
+ ua = 3.4334258940259e-09 lua = -1.5786862983809e-15
+ ub = 7.254333458e-19 lub = -1.80834088662702e-26
+ uc = 5.181291727e-13 luc = -9.76670899893637e-19
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0272246761687 lu0 = -7.98449229891865e-9
+ a0 = 0.997663879725999 la0 = -1.39553870113111e-7
+ keta = 0.04266318224 lketa = -1.12690999606489e-07 wketa = 1.05879118406788e-22 pketa = -1.0097419586829e-28
+ a1 = 0.0
+ a2 = 0.5
+ ags = -0.28313755697 lags = 9.18527068470665e-07 pags = -1.61558713389263e-27
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.158164876157715+0*(0.009/sqrt(l*w*mult))} lvoff = 7.1161645399112e-8
+ nfactor = {0.900662458620001+0*(0.02/sqrt(l*w*mult))} lnfactor = 7.33552479733592e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.4424975e-05 lcit = -8.341055750125e-12
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.271025005895605 leta0 = -2.39818499988167e-7
+ etab = -0.02847850446 letab = 2.52033340545777e-8
+ dsub = 0.0710074050500005 ldsub = 4.18737680767776e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.0769756203084007 lpclm = 9.96625507842668e-7
+ pdiblc1 = 0.00331213796900021 lpdiblc1 = 3.50647640826125e-7
+ pdiblc2 = 0.0058837902087835 lpdiblc2 = -3.87415898724586e-9
+ pdiblcb = -0.401999 lpdiblcb = 3.33642230005e-7
+ drout = 1.52153692559705 ldrout = -9.83094497065811e-7
+ pscbe1 = 429292893.4686 lpscbe1 = -114.883496156744
+ pscbe2 = 1.453303481712e-08 lpscbe2 = 1.90576441778914e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -6.0014119919695e-05 lalpha0 = 1.13126504477526e-10 walpha0 = 2.7954863898317e-26 palpha0 = -9.20368818501741e-32
+ alpha1 = 1.884995e-10 lalpha1 = -1.668211150025e-16
+ beta0 = -38.730102860375 lbeta0 = 7.86610352412926e-05 pbeta0 = -2.58493941422821e-26
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 6.146987834e-09 lagidl = 1.94646876984917e-15
+ bgidl = 805214344.000001 lbgidl = 782.057387131721
+ cgidl = 557.536247250001 lcgidl = -0.000167738631135014
+ egidl = 3.0805973382958 legidl = -2.03692057970089e-6
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.507475325 lkt1 = -1.08433724751625e-7
+ kt2 = -0.019032
+ at = 257707.396 lat = -0.20151990692302
+ ute = -1.346192304 lute = -1.01427237921522e-7
+ ua1 = 5.524e-10
+ ub1 = -3.726242641e-18 lub1 = 1.19777560571797e-25
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.81e-6
+ sbref = 2.81e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.29 pmos
* DC IV MOS Parameters
+ lmin = 8.0e-07 lmax = 1e-06 wmin = 7e-06 wmax = 1.0e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.973414853525004+0*(0.0/sqrt(l*w*mult))} lvth0 = 2.68523886603564e-8
+ k1 = 0.589870423500002 lk1 = -9.27512239538251e-9
+ k2 = 0.0154175197875001 lk2 = 1.30079044966614e-8
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 6575.92405749997 lvsat = 0.0365618656437328
+ ua = -7.35595979759993e-10 lua = 2.11087721481025e-15
+ ub = 3.83679714e-18 lub = -2.7716248099143e-24 pub = 5.60519385729927e-45
+ uc = 5.8546574915e-12 luc = -5.69947177939004e-18 wuc = -1.23259516440783e-32
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0152595189825001 lu0 = 2.60461198508241e-9
+ a0 = 0.827867713375003 la0 = 1.07148881266894e-8
+ keta = -0.15139736295 lketa = 5.90516125839353e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.869940759200002 lags = -1.01941475948204e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0946561577387+0*(0.009/sqrt(l*w*mult))} lvoff = 1.49567471418758e-8
+ nfactor = {1.54037863075+0*(0.02/sqrt(l*w*mult))} lnfactor = 1.67406865979401e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -1.2124875e-05 lcit = 1.5155428750625e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -8.59460481489988e-06 leta0 = 4.48812867021008e-11
+ etab = 0.00072873193075 letab = -6.44924115054096e-10
+ dsub = 1.4666427665 ldsub = -8.16392635938668e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.99395583862875 lpclm = -6.99892400469749e-7
+ pdiblc1 = 0.202826969022751 lpdiblc1 = 1.74078012917712e-7
+ pdiblc2 = -0.0324173066339675 lpdiblc2 = 3.00221202131046e-08 wpdiblc2 = -2.64697796016969e-23 ppdiblc2 = 1.26217744835362e-29
+ pdiblcb = -0.025
+ drout = 0.338402093148501 ldrout = 6.39739139769935e-8
+ pscbe1 = -44797159.5074997 lpscbe1 = 304.68383027684
+ pscbe2 = 1.815406017615e-08 lpscbe2 = -3.18553169343687e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.00024102438742525 lalpha0 = -1.53291069330214e-10
+ alpha1 = 0.0
+ beta0 = 66.6140227201249 lbeta0 = -1.4567989176822e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -1.97510465999997e-09 lagidl = 9.13448001657672e-15
+ bgidl = 1283382960 lbgidl = 358.8805528148
+ cgidl = -152.596199999999 lcgidl = 0.000460725034019
+ egidl = 1.79942371219525 legidl = -9.03088326470034e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.583762837500002 lkt1 = -4.09196576266879e-8
+ kt2 = -0.019032
+ at = 47124.8750000001 lat = -0.015155428750625
+ ute = -1.395725475 lute = -5.75906292523759e-8
+ ua1 = 5.524e-10
+ ub1 = -3.5909e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.41e-6
+ sbref = 2.41e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.30 pmos
* DC IV MOS Parameters
+ lmin = 6e-07 lmax = 8.0e-07 wmin = 7e-06 wmax = 1.0e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.881892254404999+0*(0.0/sqrt(l*w*mult))} lvth0 = -3.58401341238471e-8
+ k1 = 0.59352307275 lk1 = -1.17771688683865e-8
+ k2 = 0.0189560867925 lk2 = 1.05840037910715e-8
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 61502.5565075 lvsat = -0.00106260295135496
+ ua = -1.8233767778005e-09 lua = 2.85600162256401e-15
+ ub = 2.469434477865e-18 lub = -1.83498822316514e-24 wub = 2.93873587705572e-39 pub = 1.40129846432482e-45
+ uc = 2.53255847e-12 luc = -3.42385056015765e-18
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.00709052591749998 lu0 = 8.20033138964208e-9
+ a0 = 0.934519311749998 la0 = -6.23409235021911e-8
+ keta = 0.011718082125 lketa = -5.26816517152144e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = -0.561400778000001 lags = 8.78520320326111e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {0.00731538466477488+0*(0.009/sqrt(l*w*mult))} lvoff = -5.48932495467926e-8
+ nfactor = {1.78668573025+0*(0.02/sqrt(l*w*mult))} lnfactor = -1.31226564259923e-9
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -0.0573036120981399 leta0 = 3.92916817945423e-08 weta0 = 7.03103520670074e-23 peta0 = 2.52435489670724e-29
+ etab = -0.00072873193075 letab = 3.53431342754096e-10
+ dsub = 0.1933921039715 ldsub = 5.57777016400423e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.25744420752125 lpclm = 4.89609384280732e-7
+ pdiblc1 = 0.189717426328751 lpdiblc1 = 1.83057984115388e-7
+ pdiblc2 = 0.02598707339889 lpdiblc2 = -9.98458808750267e-9
+ pdiblcb = -0.025
+ drout = -0.682593035841499 ldrout = 7.63350472359498e-7
+ pscbe1 = 430689610.609 lpscbe1 = -21.022229819112
+ pscbe2 = 1.0686514267575e-08 lpscbe2 = 1.92969991620746e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -0.000115023676316125 lalpha0 = 9.06000740923091e-11 walpha0 = 2.06795153138257e-25
+ alpha1 = 0.0
+ beta0 = 27.3652154283499 lbeta0 = 1.23172475740073e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 2.30942115275e-08 lagidl = -8.03787622527987e-15
+ bgidl = 2050039997.5 lbgidl = -166.275684587514
+ cgidl = 1223.24275 lcgidl = -0.00048171776753625
+ egidl = -0.21208199437 legidl = 4.74783024998628e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.7041728745 lkt1 = 4.15606156681274e-8
+ kt2 = -0.019032
+ at = 41974.825 lat = -0.011627670250875
+ ute = -1.6071111875 lute = 8.72075268815633e-8
+ ua1 = 5.5336999e-10 lua1 = -6.64438300049995e-19
+ ub1 = -4.2982652075e-18 lub1 = 4.8454163031146e-25
+ uc1 = -2.733805074e-10 luc1 = 1.12462826666463e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.02e-6
+ sbref = 2.01e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.31 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 6e-07 wmin = 7e-06 wmax = 1.0e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.02/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.852324305450574+0*(0.0/sqrt(l*w*mult))} lvth0 = -5.01804415269973e-08 wvth0 = -5.17907185965829e-07 pvth0 = 2.51182395657492e-13
+ k1 = 0.458361440000001 lk1 = 5.37755472072001e-8
+ k2 = 0.0397051464285314 lk2 = 5.20813612894451e-10 wk2 = -1.85976049486569e-08 pk2 = 9.01974541207338e-15
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 17998.2521298435 lvsat = 0.0200367671502866 wvsat = 0.154405260891687 pvsat = -7.48857795061637e-8
+ ua = 1.1418948593867e-08 lua = -3.5664599710679e-15 wua = -8.04129742903095e-17 pua = 3.89998904659636e-23
+ ub = -5.8595928997914e-18 lub = 2.20454840986133e-24 wub = -9.67887974051201e-24 pub = 4.69420827974963e-30
+ uc = -1.62221272500001e-12 luc = -1.40880730443863e-18
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.034368285477701 lu0 = -5.02924560825759e-09 wu0 = 5.47365431085949e-08 pu0 = -2.65469497249529e-14
+ a0 = 0.214396682999999 la0 = 2.86914950828414e-7
+ keta = -0.13938919825 lketa = 2.06046237302587e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 1.25
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1225417579515+0*(0.009/sqrt(l*w*mult))} lvoff = 8.08681533638781e-9
+ nfactor = {0.704070049933691+0*(0.02/sqrt(l*w*mult))} lnfactor = 5.2375092623241e-07 wnfactor = 2.86096165448023e-06 pnfactor = -1.38755209761464e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 2.924975e-05 lcit = -9.33603250125e-12
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.0126821782940209 leta0 = 5.34892338329621e-09 weta0 = -1.44546724676185e-06 peta0 = 7.01044387343263e-13
+ etab = 0.0593853377594411 letab = -2.88015918866401e-08 wetab = -3.1284602149796e-07 petab = 1.51728756196403e-13
+ dsub = 0.419003534557 ldsub = -5.3642714136772e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.37380733260392 lpclm = -5.36816149568739e-07 wpclm = -9.65379102975844e-06 ppclm = 4.6820403804777e-12
+ pdiblc1 = 1.618697765494 lpdiblc1 = -5.09990335478063e-7
+ pdiblc2 = 0.00770696779004999 lpdiblc2 = -1.11882826774331e-9
+ pdiblcb = -0.025
+ drout = 0.859530092143 ldrout = 1.5428465902656e-8
+ pscbe1 = 482455064.78 lpscbe1 = -46.1282162647763
+ pscbe2 = 1.53528728706e-08 lpscbe2 = -3.33460674466663e-16
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -2.58245787588002e-05 lalpha0 = 4.73389577724943e-11
+ alpha1 = 0.0
+ beta0 = 45.35976918235 lbeta0 = 3.58997897608615e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 2.707805201313e-08 lagidl = -9.970018941608e-15 wagidl = -2.43755016317344e-13 pagidl = 1.1821996413883e-19
+ bgidl = 2284692500.0 lbgidl = -280.080975037499
+ cgidl = -717.926441483113 lcgidl = 0.000459739584487102 wcgidl = 0.00816850143570121 pcgidl = -3.96168235380791e-9
+ egidl = 1.15799168033 legidl = -1.89695856862498e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.67622925 lkt1 = 2.80080975037504e-8
+ kt2 = -0.019032
+ at = 18000.0
+ ute = -1.638662255 lute = 1.02509636863725e-7
+ ua1 = 5.52e-10
+ ub1 = -7.68506304000001e-18 lub1 = 2.1271216450848e-24
+ uc1 = -4.1496e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 1.81e-6
+ sbref = 1.81e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.32 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.996534475654001+0*(0.0/sqrt(l*w*mult))} wvth0 = 1.22974172098248e-7
+ k1 = 0.59521
+ k2 = 0.021882733159 wk2 = -2.29100635895282e-10
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200000.0
+ ua = 2.70536302101584e-09 wua = -3.78685728008627e-18
+ ub = 1.4287104508e-19 wub = -1.12012587826951e-24
+ uc = -3.9972e-11
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0226695689992 wu0 = -9.06533593111757e-9
+ a0 = 0.8913783700167 wa0 = 1.08047384513407e-8
+ keta = -0.0079259
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.151862771388 wags = -4.43397846086551e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.093204657+0*(0.009/sqrt(l*w*mult))}
+ nfactor = {1.7272132821+0*(0.02/sqrt(l*w*mult))} wnfactor = 2.69633825322902e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.0800000000000101
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.08353125
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0029407877
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 333712830.0
+ pscbe2 = 1.5000958e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 5.0667189e-5
+ alpha1 = 0.0
+ beta0 = 38.266046
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -1.27169970729e-08 wagidl = 1.40990293642535e-13
+ bgidl = 1704700000.0
+ cgidl = -53.0729000000001 wcgidl = 0.0052869377514294
+ egidl = 0.69350825
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.57505223439 wkt1 = -4.7582439762857e-9
+ kt2 = -0.019032
+ at = 382807.4316 wat = 0.331314765756243
+ ute = -1.0106166229 wute = -2.63818193796326e-6
+ ua1 = 2.424730964752e-09 wua1 = -1.20623952036479e-14
+ ub1 = -1.8454471989e-18 wub1 = -9.12349224638334e-24
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.33 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.996534475653999+0*(0.0/sqrt(l*w*mult))} wvth0 = 1.22974172098251e-7
+ k1 = 0.59521
+ k2 = 0.021882733159 wk2 = -2.29100635895176e-10
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200000.0
+ ua = 2.70536302101584e-09 wua = -3.78685728008627e-18
+ ub = 1.4287104508e-19 wub = -1.12012587826951e-24
+ uc = -3.9972e-11
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0226695689992 wu0 = -9.06533593111757e-9
+ a0 = 0.8913783700167 wa0 = 1.08047384513407e-8
+ keta = -0.0079259
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.151862771388 wags = -4.43397846086559e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.093204657+0*(0.009/sqrt(l*w*mult))}
+ nfactor = {1.7272132821+0*(0.02/sqrt(l*w*mult))} wnfactor = 2.69633825322902e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.0800000000000101
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.08353125
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0029407877
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 333712830.0
+ pscbe2 = 1.5000958e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 5.0667189e-5
+ alpha1 = 0.0
+ beta0 = 38.266046
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -1.27169970729e-08 wagidl = 1.40990293642536e-13
+ bgidl = 1704700000.0
+ cgidl = -53.0728999999997 wcgidl = 0.00528693775142941
+ egidl = 0.69350825
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.57505223439 wkt1 = -4.75824397628232e-9
+ kt2 = -0.019032
+ at = 382807.4316 wat = 0.331314765756243
+ ute = -1.0106166229 wute = -2.63818193796327e-6
+ ua1 = 2.424730964752e-09 wua1 = -1.20623952036479e-14
+ ub1 = -1.8454471989e-18 wub1 = -9.12349224638333e-24
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.34 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.00077795304219+0*(0.0/sqrt(l*w*mult))} lvth0 = 3.34597979885031e-08 wvth0 = 1.10598986743659e-07 pvth0 = 9.75782746450203e-14
+ k1 = 0.6040969260625 lk1 = -7.0073367568183e-8
+ k2 = 0.0204326382859806 lk2 = 1.14339908232835e-08 wk2 = -6.20958440200139e-09 pk2 = 4.71560845933275e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 357823.114873562 lvsat = -1.24443447166246 wvsat = -0.4261993296395 pvsat = 3.36057958321081e-6
+ ua = 2.45152509007856e-09 lua = 2.00151081625081e-15 wua = -8.35127384660568e-19 pua = -2.32743754668239e-23
+ ub = 3.3831329261499e-19 lub = -1.54106114460216e-24 wub = -6.90332096452327e-25 pub = -3.38892182065958e-30
+ uc = -5.150363640875e-11 luc = 9.09268954248117e-17
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0218445699958255 lu0 = 6.50511301661283e-09 wu0 = -7.94420918045944e-09 pu0 = -8.84007882330577e-15
+ a0 = 0.916242157490703 la0 = -1.96050839913581e-07 wa0 = -2.27941978822848e-08 pa0 = 2.64927444995913e-13
+ keta = -0.004975149172625 lketa = -2.32666555200977e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.104290491958294 lags = 3.75107185441838e-07 wags = 1.05687514356132e-07 pags = -1.18296450220084e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0947667260771125+0*(0.009/sqrt(l*w*mult))} lvoff = 1.23169068626865e-8
+ nfactor = {1.82091157948594+0*(0.02/sqrt(l*w*mult))} lnfactor = -7.38810606396655e-07 wnfactor = -3.35261126864248e-07 pnfactor = 4.7695936735209e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.0800000000000101
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.643778489125225 lpclm = 5.7348336564537e-06 wpclm = 4.2351647362715e-22 ppclm = 6.46234853557053e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00454411319014037 lpdiblc2 = -1.26422134731294e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 560706123.996462 lpscbe1 = -1789.84098819564
+ pscbe2 = -1.51292780647975e-08 lpscbe2 = 2.37576760719748e-13 ppscbe2 = -3.85185988877447e-34
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 7.7982685969875e-05 lalpha0 = -2.1538255702998e-10
+ alpha1 = 0.0
+ beta0 = 39.1348639430787 lbeta0 = -6.85062513708606e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -3.38140076936816e-08 lagidl = 1.6634982325981e-13 wagidl = 2.83332311522658e-13 pagidl = -1.12236609927468e-18
+ bgidl = 1298122546.492 lbgidl = 3205.86118802327 wbgidl = 1275.17470113023 pbgidl = -0.0100547461425384
+ cgidl = -70.5988758465182 lcgidl = 0.000138192231919916 wcgidl = 0.00703281452344663 pcgidl = -1.3766229617972e-8
+ egidl = 1.20611845100666 legidl = -4.04192887188653e-6
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.608224909485457 lkt1 = 2.61566377264305e-07 wkt1 = 1.61784706923003e-07 pkt1 = -1.31319033512615e-12
+ kt2 = -0.019032
+ at = 711118.207917427 lat = -2.58872882970903 wat = -0.277859296166241 pat = 4.80333443238847e-6
+ ute = -0.480816574745845 lute = -4.17747073069526e-06 wute = -5.20051284748267e-06 pute = 2.0203966409906e-11
+ ua1 = 4.75828717097368e-09 lua1 = -1.84000790182769e-14 wua1 = -2.37779814671969e-14 pua1 = 9.23773391101528e-20
+ ub1 = -5.02052890422302e-19 lub1 = -1.05926574053751e-23 wub1 = -1.48249780577455e-23 pub1 = 4.49561871151615e-29
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.35 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.977341782321512+0*(0.0/sqrt(l*w*mult))} lvth0 = -5.75896080804813e-08 wvth0 = 1.33853738874992e-07 pvth0 = 7.23367888853917e-15
+ k1 = 0.6023840567 lk1 = -6.34188786592171e-8
+ k2 = 0.0216365998351186 lk2 = 6.7566062246898e-09 wk2 = 1.82711262762731e-08 pk2 = -4.7951353988215e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -13015.3867031982 lvsat = 0.196271252770746 wvsat = 0.686301138833073 pvsat = -9.61479174302793e-7
+ ua = 3.3160868828489e-09 lua = -1.35730742585302e-15 wua = -1.25734378308553e-17 pua = 2.23289019251281e-23
+ ub = -8.28255519361864e-19 lub = 2.99105285708386e-24 wub = -2.75306349710012e-24 pub = 4.62477935720008e-30
+ uc = -5.45822372525e-11 luc = 1.02887244309776e-16
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0229736663168666 lu0 = 2.11857945484981e-09 wu0 = -1.25154506011168e-08 pu0 = 8.91917123974039e-15
+ a0 = 0.813514281650165 la0 = 2.0304644408753e-07 wa0 = 7.23170929937135e-08 pa0 = -1.04579444500868e-13
+ keta = -0.00516198539000001 lketa = -2.2540797749777e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.180805358651186 lags = 7.78473109142846e-08 wags = -2.67361674505817e-07 pags = 2.66329731281876e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0644364973897326+0*(0.009/sqrt(l*w*mult))} lvoff = -1.05515879936641e-7
+ nfactor = {1.73956705973018+0*(0.02/sqrt(l*w*mult))} lnfactor = -4.22787553868146e-07 wnfactor = 3.2253744256166e-06 pnfactor = -9.06345764468949e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.01986865950001 leta0 = 2.33609957185798e-7
+ etab = -0.12173557277 letab = 2.00992441533586e-7
+ dsub = 0.811505457874999 ldsub = -9.77097446317086e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.04601663892438 lpclm = -8.30011967043352e-7
+ pdiblc1 = 0.5791285228315 lpdiblc1 = -7.34763365557764e-7
+ pdiblc2 = -0.00110255629368 lpdiblc2 = 9.29506923816533e-9
+ pdiblcb = 0.1634995 lpdiblcb = -7.323196150025e-07 ppdiblcb = 6.05845175209737e-28
+ drout = 0.1453011 ldrout = 1.6111031530055e-6
+ pscbe1 = -152915980.78355 lpscbe1 = 982.577320764188 ppscbe1 = 8.67361737988404e-19
+ pscbe2 = 7.56929177375625e-08 lpscbe2 = -1.15267015861442e-13 wpscbe2 = 2.01948391736579e-28
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 4.37897997750275e-05 lalpha0 = -8.2543365127428e-11
+ alpha1 = -9.424975e-11 lalpha1 = 3.6615980750125e-16
+ beta0 = 69.7665703037275 lbeta0 = -0.000125854651189675
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.66927448378717e-08 lagidl = -2.9868657791512e-14 wagidl = -5.27105033430435e-14 pagidl = 1.831585562645e-19
+ bgidl = 2974589195.51599 lbgidl = -3307.20336110167 wbgidl = -2550.34940226047 pbgidl = 0.00480739587151396
+ cgidl = -509.649227499716 lcgidl = 0.00184390065284083 wcgidl = 0.00677810982077278 pcgidl = -1.27767031216076e-8
+ egidl = -1.56307736015895 legidl = 6.71638300851282e-06 wegidl = -8.470329472543e-22 pegidl = 9.69352280335579e-27
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.5418400675 lkt1 = 3.6615980750127e-09 wkt1 = -1.76231258380978e-7
+ kt2 = -0.019032
+ at = -163978.993357488 lat = 0.811019421758009 wat = 2.62597482209082 pat = -6.47804659786962e-6
+ ute = -1.82104556779425 lute = 1.02931220615281e-06 wute = 8.27165651820722e-07 pute = -3.21353442149524e-12
+ ua1 = -4.7771419424e-10 lua1 = 1.94176010557143e-15 wua1 = -9.86076131526265e-32 pua1 = 3.76158192263132e-37
+ ub1 = -2.64960813536477e-18 lub1 = -2.24941601654986e-24 wub1 = -7.51196945394647e-24 pub1 = 1.65451852544454e-29
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.36 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.09122170905861+0*(0.0/sqrt(l*w*mult))} lvth0 = 1.57073484419306e-07 wvth0 = 4.41817501106195e-07 pvth0 = -5.73276473098463e-13
+ k1 = 0.55931480325 lk1 = 1.77664487477661e-8
+ k2 = 0.0147963264130086 lk2 = 1.96504874240002e-08 wk2 = 2.92642546783611e-08 pk2 = -6.86733460605089e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 129355.78835715 lvsat = -0.0720977003621359 wvsat = 0.332195040891855 pvsat = -2.93990950214088e-7
+ ua = 3.43512544151842e-09 lua = -1.58169451375226e-15 wua = -1.19316493775657e-17 pua = 2.1119133899577e-23
+ ub = 1.94992897776354e-18 lub = -2.24581102907505e-24 wub = -8.59655444126122e-24 pub = 1.5639730569489e-29
+ uc = 5.181291727e-13 luc = -9.76670899893637e-19
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.031774629556353 lu0 = -1.4471192246766e-08 wu0 = -3.19428840586708e-08 pu0 = 4.55397861700627e-14
+ a0 = 1.00080303533473 la0 = -1.49991920164113e-07 wa0 = -2.20383980029448e-08 pa0 = 7.32801842503644e-14
+ keta = 0.04266318224 lketa = -1.12690999606489e-7
+ a1 = 0.0
+ a2 = 0.5
+ ags = -0.23772850061783 lags = 8.66781542967083e-07 wags = -3.18793644393625e-07 pags = 3.63278737360549e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.208611890413665+0*(0.009/sqrt(l*w*mult))} lvoff = 1.66254015036506e-07 wvoff = 3.54162557325696e-07 pvoff = -6.67594649746151e-13
+ nfactor = {0.903513996818727+0*(0.02/sqrt(l*w*mult))} lnfactor = 1.15316828945463e-06 wnfactor = -2.00191840026427e-08 pnfactor = -2.94590691752525e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.4424975e-05 lcit = -8.34105575012501e-12
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.272101061503416 leta0 = -2.41846859428613e-07 weta0 = -7.55443332985742e-09 peta0 = 1.42400690546153e-14
+ etab = -0.02847850446 letab = 2.52033340545777e-8
+ dsub = -0.473650622302969 ldsub = 1.44541533903798e-06 wdsub = 3.82376405581914e-06 pdsub = -7.20777612639879e-12
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.0769756203083998 lpclm = 9.96625507842668e-7
+ pdiblc1 = 0.00331213796900021 lpdiblc1 = 3.50647640826125e-7
+ pdiblc2 = 0.0058837902087835 lpdiblc2 = -3.87415898724585e-9
+ pdiblcb = -0.401999 lpdiblcb = 3.33642230005e-07 ppdiblcb = 8.07793566946316e-28
+ drout = 1.52153692559705 ldrout = -9.83094497065812e-7
+ pscbe1 = 429292893.4686 lpscbe1 = -114.883496156744
+ pscbe2 = 1.453303481712e-08 lpscbe2 = 1.90576441778787e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -6.0014119919695e-05 lalpha0 = 1.13126504477526e-10 walpha0 = -5.87448938899983e-26 palpha0 = 4.38562836359586e-33
+ alpha1 = 1.884995e-10 lalpha1 = -1.668211150025e-16
+ beta0 = -38.730102860375 lbeta0 = 7.86610352412926e-05 pbeta0 = -5.16987882845642e-26
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -3.72917171183784e-09 lagidl = 8.62655279510771e-15 wagidl = 6.9335439825321e-14 pagidl = -4.68974363781513e-20
+ bgidl = 527298125.776496 lbgidl = 1305.92806890193 wbgidl = 1951.10691921105 pbgidl = -0.00367782678717824
+ cgidl = 557.53624725 lcgidl = -0.000167738631135013 wcgidl = 1.73472347597681e-18
+ egidl = 3.0805973382958 legidl = -2.03692057970089e-6
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.46015736996215 lkt1 = -1.50309878370347e-07 wkt1 = -3.32195040891853e-07 pkt1 = 2.93990950214086e-13
+ kt2 = -0.019032
+ at = 475369.98917411 lat = -0.394150213569142 wat = -1.52809718810254 pat = 1.3523583709848e-6
+ ute = -1.11054888791151 lute = -3.09970482942757e-07 wute = -1.65433130364144e-06 pute = 1.46407493206616e-12
+ ua1 = 5.524e-10
+ ub1 = -4.06598555817176e-18 lub1 = 4.20448343554217e-25 wub1 = 2.38516039360353e-24 pub1 = -2.11085502253715e-30
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.81e-6
+ sbref = 2.81e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.37 pmos
* DC IV MOS Parameters
+ lmin = 8.0e-07 lmax = 1e-06 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.775578190861344+0*(0.0/sqrt(l*w*mult))} lvth0 = -1.22269450967681e-07 wvth0 = -1.38890952051692e-06 pvth0 = 1.04690778740288e-12
+ k1 = 0.589870423500001 lk1 = -9.27512239538251e-9
+ k2 = 0.0412132161731274 lk2 = -3.72832792925614e-09 wk2 = -1.81098325335547e-07 pk2 = 1.174964854389e-13
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 3604.62131175934 lvsat = 0.0391914537171993 wvsat = 0.0208599893282329 pvsat = -1.84609862555393e-8
+ ua = -7.50524998045325e-10 lua = 2.12258519700946e-15 wua = 1.0480896386586e-16 pua = -8.21957251177961e-23
+ ub = -2.05018430546795e-18 lub = 1.29426922601841e-24 wub = 4.13294708201675e-23 pub = -2.85445521567491e-29
+ uc = 5.8546574915e-12 luc = -5.69947177939004e-18 puc = 5.87747175411144e-39
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.00150216967633571 lu0 = 1.23197833847499e-08 wu0 = 9.65832782010356e-08 pu0 = -6.82052247989661e-14
+ a0 = 0.789568148209744 la0 = 3.69498987670637e-08 wa0 = 2.68881561048747e-07 pa0 = -1.84182524910583e-13
+ keta = -0.15139736295 lketa = 5.90516125839353e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.812147070814031 lags = -6.2353088372258e-08 wags = 4.05739780202043e-07 pags = -2.779297207395e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {0.157578913541049+0*(0.009/sqrt(l*w*mult))} lvoff = -1.57823015509396e-07 wvoff = -1.77081278662848e-06 pvoff = 1.21299790477657e-12
+ nfactor = {3.42478895085802+0*(0.02/sqrt(l*w*mult))} lnfactor = -1.07814743849537e-06 wnfactor = -1.32294762705739e-05 pnfactor = 8.7443965568049e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -1.2124875e-05 lcit = 1.5155428750625e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.00023944192407801 leta0 = -1.25068540899633e-09 weta0 = -1.7413369785813e-09 peta0 = 9.09550784921709e-15
+ etab = -0.00201516642371491 letab = 1.78341220915558e-09 wetab = 1.9263499982944e-08 petab = -1.70481011674055e-14
+ dsub = 4.18996308055835 ldsub = -2.68185946992577e-06 wdsub = -1.91190321383623e-05 pdsub = 1.30964837914708e-11
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.99395583862875 lpclm = -6.9989240046975e-7
+ pdiblc1 = 0.202826969022749 lpdiblc1 = 1.74078012917711e-7
+ pdiblc2 = -0.0324173066339675 lpdiblc2 = 3.00221202131046e-08 wpdiblc2 = -1.32348898008484e-23 ppdiblc2 = -3.78653234506086e-29
+ pdiblcb = -0.025
+ drout = 0.3384020931485 ldrout = 6.39739139769935e-8
+ pscbe1 = -44797159.5075006 lpscbe1 = 304.683830276841
+ pscbe2 = 1.815406017615e-08 lpscbe2 = -3.18553169343687e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.00024102438742525 lalpha0 = -1.53291069330214e-10
+ alpha1 = 0.0
+ beta0 = 66.6140227201249 lbeta0 = -1.45679891768221e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 3.3685895728122e-08 lagidl = -2.44855948139195e-14 wagidl = -2.50357553970805e-13 pagidl = 2.36029264666451e-19
+ bgidl = 2672964051.11752 lbgidl = -592.975546695241 wbgidl = -9755.53459605527 pbgidl = 0.00668249242062487
+ cgidl = -152.5962 lcgidl = 0.000460725034019001
+ egidl = 1.79942371219525 legidl = -9.03088326470035e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.557970278943223 lkt1 = -6.374594298664e-08 wkt1 = -1.81076296252021e-07 pkt1 = 1.60251616801556e-13
+ kt2 = -0.019032
+ at = 47124.8749999999 lat = -0.015155428750625
+ ute = -1.395725475 lute = -5.75906292523742e-8
+ ua1 = 5.524e-10
+ ub1 = -3.5909e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.41e-6
+ sbref = 2.41e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.38 pmos
* DC IV MOS Parameters
+ lmin = 6e-07 lmax = 8.0e-07 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.949915828838735+0*(0.0/sqrt(l*w*mult))} lvth0 = -2.84904064135833e-09 wvth0 = 4.77558551981999e-07 pvth0 = -2.31613509918506e-13
+ k1 = 0.59352307275 lk1 = -1.17771688683865e-8
+ k2 = 0.0236245398912763 lk2 = 8.31982738043044e-09 wk2 = -3.27748096216158e-08 pk2 = 1.58956187924355e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 64473.8592532405 lvsat = -0.0025036699265254 wvsat = -0.0208599893282329 pvsat = 1.01169905242462e-8
+ ua = -1.81596838120624e-09 lua = 2.85240858725778e-15 wua = -5.20105445724568e-17 pua = 2.52248540649256e-23
+ ub = 2.63614038133696e-18 lub = -1.91583975281952e-24 wub = -1.17035646144222e-24 pub = 5.67617032017169e-31
+ uc = 2.53255847000001e-12 luc = -3.42385056015765e-18
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.00854780547595779 lu0 = 7.49355809018786e-09 wu0 = -1.02308107382391e-08 pu0 = 4.96189205399226e-15
+ a0 = 0.93451931175 la0 = -6.23409235021911e-8
+ keta = 0.0117180821250001 lketa = -5.26816517152144e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = -0.561400777999999 lags = 8.7852032032611e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {0.00731538466477499+0*(0.009/sqrt(l*w*mult))} lvoff = -5.48932495467926e-8
+ nfactor = {2.0129724439881+0*(0.02/sqrt(l*w*mult))} lnfactor = -1.11060190372012e-07 wnfactor = -1.58864270578437e-06 pnfactor = 7.70483769091895e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -0.062931926666087 leta0 = 4.20213862184238e-08 weta0 = 3.95135036278689e-08 peta0 = -1.91638516919983e-14
+ etab = 0.00201516642371492 letab = -9.77345639669616e-10 wetab = -1.9263499982944e-08 petab = 9.34270117422791e-15
+ dsub = 0.193361926677988 ldsub = 5.5792337476509e-08 wdsub = 2.11859266614149e-10 pdsub = -1.02750685011713e-16
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.25744420752125 lpclm = 4.89609384280732e-7
+ pdiblc1 = 0.18971742632875 lpdiblc1 = 1.83057984115388e-7
+ pdiblc2 = 0.02598707339889 lpdiblc2 = -9.98458808750267e-9
+ pdiblcb = -0.025
+ drout = -0.682593035841501 ldrout = 7.63350472359499e-7
+ pscbe1 = 430689610.609 lpscbe1 = -21.022229819112
+ pscbe2 = 1.0686514267575e-08 lpscbe2 = 1.92969991620746e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -0.000115023676316125 lalpha0 = 9.0600074092309e-11 walpha0 = -2.06795153138257e-25 palpha0 = 9.86076131526265e-32
+ alpha1 = 0.0
+ beta0 = 27.36521542835 lbeta0 = 1.23172475740074e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -2.28681278206731e-08 lagidl = 1.42536285468873e-14 wagidl = 3.22677959921098e-13 pagidl = -1.56497197171933e-19
+ bgidl = 2050039997.5 lbgidl = -166.27568458751
+ cgidl = 1223.24275 lcgidl = -0.00048171776753625
+ egidl = -0.212081994370001 legidl = 4.74783024998628e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.729965433056775 lkt1 = 5.40698776053706e-08 wkt1 = 1.81076296252021e-07 pkt1 = -8.7821098300747e-14
+ kt2 = -0.019032
+ at = 41974.825 lat = -0.011627670250875
+ ute = -1.6071111875 lute = 8.72075268815616e-8
+ ua1 = 5.53369989999999e-10 lua1 = -6.64438300049995e-19
+ ub1 = -4.2982652075e-18 lub1 = 4.8454163031146e-25
+ uc1 = -2.733805074e-10 luc1 = 1.12462826666463e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.02e-6
+ sbref = 2.01e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.39 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 6e-07 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.07881637645913+0*(0.0/sqrt(l*w*mult))} lvth0 = 5.96670804517951e-08 wvth0 = 1.07217722766072e-06 pvth0 = -5.20000594529314e-13
+ k1 = 0.345578941858291 lk1 = 1.08474494893439e-07 wk1 = 7.91787949248905e-07 pk1 = -3.8401319644597e-13
+ k2 = 0.0277590320935883 lk2 = 6.31461933477017e-09 wk2 = 6.52699234942106e-08 pk2 = -3.16555865450747e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 98401.9043477615 lvsat = -0.0189586021571427 wvsat = -0.410067453853078 pvsat = 1.98880664781474e-7
+ ua = 1.78992016965993e-08 lua = -6.70935032462753e-15 wua = -4.55749391584788e-14 pua = 2.21036176171664e-20
+ ub = -7.56152642249609e-18 lub = 3.02997765870549e-24 wub = 2.26952072856691e-24 pub = -1.1007062057513e-30
+ uc = -4.57513852198308e-11 luc = 1.99936207096918e-17 wuc = 3.09808237691544e-16 puc = -1.50255446239211e-22
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0675308886263449 lu0 = -2.11129423223342e-08 wu0 = -1.78081048020016e-07 pu0 = 8.63684178844676e-14
+ a0 = -1.33972101418666 la0 = 1.04065426337546e-06 wa0 = 1.09106615354512e-05 pa0 = -5.29161629138615e-12
+ keta = -0.0405619638029457 lketa = -2.73260908403903e-08 wketa = -6.93815215854262e-07 pketa = 3.36496910613238e-13
+ a1 = 0.0
+ a2 = 0.5
+ ags = 1.25
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.426185681461714+0*(0.009/sqrt(l*w*mult))} lvoff = 1.55352600019224e-07 wvoff = 2.13172791398852e-06 pvoff = -1.03387737964486e-12
+ nfactor = {-5.02940629485104+0*(0.02/sqrt(l*w*mult))} lnfactor = 3.30445828607128e-06 wnfactor = 4.31127520643726e-05 pnfactor = -2.09094691874604e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 2.924975e-05 lcit = -9.33603250125e-12 wcit = 1.03397576569128e-25
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -0.577154291983696 leta0 = 2.91416662285637e-07 weta0 = 2.69547143511227e-06 peta0 = -1.30729016867228e-12
+ etab = -0.0468222719534339 letab = 2.27085677860557e-08 wetab = 4.32783015584743e-07 petab = -2.09897598643523e-13
+ dsub = 0.523562188072002 ldsub = -1.0435313829828e-07 wdsub = -7.3405256318092e-07 pdsub = 3.56011822879931e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.474509764920867 lpclm = 8.44603401145294e-07 wpclm = 1.03427792769749e-05 ppclm = -5.01619623543645e-12
+ pdiblc1 = 2.57219637615875 lpdiblc1 = -9.72432394157414e-07 wpdiblc1 = -6.69402364719134e-06 ppdiblc1 = 3.24656799876957e-12
+ pdiblc2 = 0.0383269308871603 lpdiblc2 = -1.59693572700263e-08 wpdiblc2 = -2.14967022243779e-07 ppdiblc2 = 1.04257930953122e-13
+ pdiblcb = -0.025
+ drout = -0.850467997156063 ldrout = 8.44768989222255e-07 wdrout = 1.20050176459508e-05 pdrout = -5.82237353319792e-12
+ pscbe1 = 47009764.1890898 lpscbe1 = 165.060577295313 wpscbe1 = 3057.03763656427 ppscbe1 = -0.00148264796854549
+ pscbe2 = 1.50871333374893e-08 lpscbe2 = -2.0457832960561e-16 wpscbe2 = 1.86562067185052e-15 ppscbe2 = -9.04816697744187e-22
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -0.000538554158683642 lalpha0 = 2.96010240388143e-10 walpha0 = 3.59961083764823e-09 palpha0 = -1.74579325820521e-15
+ alpha1 = 0.0
+ beta0 = 5.24832097093451 lbeta0 = 2.30438308013816e-05 wbeta0 = 0.000281601860607967 pbeta0 = -1.36575494385561e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 6.21613953927692e-09 lagidl = 1.47904298648397e-16 wagidl = -9.72942518614328e-14 pagidl = 4.71872256815356e-20
+ bgidl = 3392222430.33761 lbgidl = -817.22745360159 wbgidl = -7775.39837051617 pbgidl = 0.00377102933270849
+ cgidl = 2629.7312685541 lcgidl = -0.0011638576665924 wcgidl = -0.0153336826504071 pcgidl = 7.43675941703421e-9
+ egidl = 1.24554762326611 legidl = -2.32160051406798e-07 wegidl = -6.14685271599764e-07 pegidl = 2.98119283299525e-13
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.482943049242998 lkt1 = -6.57347434323913e-08 wkt1 = -1.35696306640771e-06 pkt1 = 6.58120302392408e-13
+ kt2 = -0.019032
+ at = 18000.0
+ ute = -1.638662255 lute = 1.02509636863725e-7
+ ua1 = 5.52e-10
+ ub1 = -1.47786666077819e-17 lub1 = 5.5674839074412e-24 wub1 = 4.9800544537163e-23 pub1 = -2.41530150978014e-29
+ uc1 = -4.1496e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 1.81e-6
+ sbref = 1.81e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.40 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.995697956595+0*(0.0/sqrt(l*w*mult))} wvth0 = 1.18774439873805e-7
+ k1 = 0.59521
+ k2 = 0.0219550499783 wk2 = -5.92166214755466e-10
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200000.0
+ ua = 2.70497525936343e-09 wua = -1.84010533281334e-18
+ ub = 4.52993958999999e-21 wub = -4.25586294932441e-25
+ uc = -3.9972e-11
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.02180956885931 wu0 = -4.74771726880185e-9
+ a0 = 0.8913176919564 wa0 = 1.1109371803581e-8
+ keta = -0.0079259
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.1558621755523 wags = -6.44187372238643e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.093204657+0*(0.009/sqrt(l*w*mult))}
+ nfactor = {1.78761037649+0*(0.02/sqrt(l*w*mult))} wnfactor = -3.35889415027755e-8
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.0800000000000101
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.08353125
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0029407877
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 333712830.0
+ pscbe2 = 1.5000958e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 5.0667189e-5
+ alpha1 = 0.0
+ beta0 = 38.266046
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.6258553613e-08 wagidl = -4.48105291831594e-15
+ bgidl = 1597472747 wbgidl = 538.332922504957
+ cgidl = 1000.0
+ egidl = 0.69350825
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.576
+ kt2 = -0.019032
+ at = 448800.0
+ ute = -1.5361
+ ua1 = 2.2096e-11
+ ub1 = -3.6627e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.41 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.995697956595+0*(0.0/sqrt(l*w*mult))} wvth0 = 1.18774439873805e-7
+ k1 = 0.59521
+ k2 = 0.0219550499783 wk2 = -5.92166214755413e-10
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200000.0
+ ua = 2.70497525936343e-09 wua = -1.84010533281334e-18
+ ub = 4.52993959000004e-21 wub = -4.25586294932441e-25
+ uc = -3.9972e-11
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.02180956885931 wu0 = -4.74771726880179e-9
+ a0 = 0.8913176919564 wa0 = 1.1109371803581e-8
+ keta = -0.0079259
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.1558621755523 wags = -6.44187372238643e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.093204657+0*(0.009/sqrt(l*w*mult))}
+ nfactor = {1.78761037649+0*(0.02/sqrt(l*w*mult))} wnfactor = -3.35889415027755e-8
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.0800000000000101
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.08353125
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0029407877
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 333712830.0
+ pscbe2 = 1.5000958e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 5.0667189e-5
+ alpha1 = 0.0
+ beta0 = 38.266046
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.6258553613e-08 wagidl = -4.48105291831592e-15
+ bgidl = 1597472747.0 wbgidl = 538.332922504957
+ cgidl = 1000.0
+ egidl = 0.69350825
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.576
+ kt2 = -0.019032
+ at = 448800.0
+ ute = -1.5361
+ ua1 = 2.2096e-11
+ ub1 = -3.6627e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.42 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.00404921193231+0*(0.0/sqrt(l*w*mult))} lvth0 = 6.58496065784092e-08 wvth0 = 1.27022296203872e-07 pvth0 = -6.50343059232972e-14
+ k1 = 0.6040969260625 lk1 = -7.0073367568183e-8
+ k2 = 0.0184917321634947 lk2 = 2.73082436531505e-08 wk2 = 3.53470761325334e-09 pk2 = -3.25403794994804e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 272931.0686375 lvsat = -0.575061111551344
+ ua = 2.45138086899304e-09 lua = 1.99959050009857e-15 wua = -1.11067443889232e-19 pua = -1.36334551089641e-23
+ ub = 3.34880065225554e-19 lub = -2.60480908888571e-24 wub = -6.73095626408846e-25 pub = 1.95160984114479e-30
+ uc = -5.150363640875e-11 luc = 9.09268954248118e-17
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0213763740588575 lu0 = 3.41573883559431e-09 wu0 = -5.59363803365442e-09 pu0 = 6.67008100125881e-15
+ a0 = 0.908628948860843 la0 = -1.36499174135248e-07 wa0 = 1.54278094590134e-08 pa0 = -3.40508593208872e-14
+ keta = -0.004975149172625 lketa = -2.32666555200977e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.142232788089719 lags = 1.07467651995514e-07 wags = -8.48012521795438e-08 pags = 1.60716028512957e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0947667260771125+0*(0.009/sqrt(l*w*mult))} lvoff = 1.23169068626867e-8
+ nfactor = {1.72693975640564+0*(0.02/sqrt(l*w*mult))} lnfactor = 4.78387536012075e-07 wnfactor = 1.36523095304868e-07 pnfactor = -1.34133255966809e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.0800000000000101
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.643778489125225 lpclm = 5.7348336564537e-06 wpclm = -4.2351647362715e-22 ppclm = -1.61558713389263e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00454411319014037 lpdiblc2 = -1.26422134731294e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 560706123.996463 lpscbe1 = -1789.84098819564
+ pscbe2 = -1.51292780647975e-08 lpscbe2 = 2.37576760719748e-13
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 7.7982685969875e-05 lalpha0 = -2.1538255702998e-10
+ alpha1 = 0.0
+ beta0 = 39.1348639430788 lbeta0 = -6.85062513708617e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 2.65867730818574e-08 lagidl = -8.14379588708432e-14 wagidl = -1.99089627500049e-14 pagidl = 1.21648991883319e-19
+ bgidl = 1340745232.93282 lbgidl = 2024.29516478218 wbgidl = 1061.18810057174 pbgidl = -0.00412271046478073
+ cgidl = 1330.224575 lcgidl = -0.00260381912275213
+ egidl = 1.20611845100666 legidl = -4.04192887188653e-6
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.576
+ kt2 = -0.019032
+ at = 646913.506004285 lat = -1.56212400427625 wat = 0.044479510922864 pat = -3.50720721229233e-7
+ ute = -1.516675025 lute = -1.53165830750129e-7
+ ua1 = 2.2096e-11
+ ub1 = -3.27453083238361e-18 lub1 = -3.06071194580939e-24 wub1 = -9.05791364819927e-25 pub1 = 7.14216038264831e-30
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.43 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.968738953469704+0*(0.0/sqrt(l*w*mult))} lvth0 = -7.13305709975179e-08 wvth0 = 9.06633570640922e-08 pvth0 = 7.6219990840051e-14
+ k1 = 0.602384056700001 lk1 = -6.34188786592171e-8
+ k2 = 0.0280785256728192 lk2 = -9.93640119660737e-09 wk2 = -1.40704722049405e-08 pk2 = 3.58556560683035e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 137918.755768925 lvsat = -0.0505389511184948 wvsat = -0.0714616103702279 pvsat = 2.77627998980282e-7
+ ua = 3.31556165379298e-09 lua = -1.35774752794527e-15 wua = -9.93653270880493e-18 pua = 2.45384283178804e-23
+ ub = -1.37278117325411e-18 lub = 4.0294462843016e-24 wub = -1.92800750932322e-26 pub = -5.88460306638609e-31
+ uc = -5.45822372525e-11 luc = 1.02887244309776e-16
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0207514137085906 lu0 = 5.84370667157918e-09 wu0 = -1.35866249280379e-09 pu0 = -9.78277780006824e-15
+ a0 = 0.827346419450145 la0 = 1.79283046212663e-07 wa0 = 2.87303881884309e-09 pa0 = 1.47243618423186e-14
+ keta = -0.00516198539000001 lketa = -2.25407977497769e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.131234105358444 lags = 1.50197479413102e-07 wags = -1.84898913471524e-08 pags = -9.69032767640774e-14
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0644364973897325+0*(0.009/sqrt(l*w*mult))} lvoff = -1.05515879936641e-7
+ nfactor = {2.60127119538399+0*(0.02/sqrt(l*w*mult))} lnfactor = -2.91838573276163e-06 wnfactor = -1.10079912357543e-06 pnfactor = 3.46565807407078e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.0198686595000102 leta0 = 2.33609957185797e-7
+ etab = -0.12173557277 letab = 2.00992441533586e-7
+ dsub = 0.811505457875 ldsub = -9.77097446317086e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.04601547173617 lpclm = -8.30007432523007e-07 wpclm = 5.85985205095398e-12 ppclm = -2.27654959187431e-17
+ pdiblc1 = 0.5791285228315 lpdiblc1 = -7.34763365557763e-7
+ pdiblc2 = -0.00110255629368 lpdiblc2 = 9.29506923816533e-9
+ pdiblcb = 0.1634995 lpdiblcb = -7.323196150025e-07 ppdiblcb = -1.0097419586829e-28
+ drout = 0.1453011 ldrout = 1.6111031530055e-6
+ pscbe1 = -152915980.78355 lpscbe1 = 982.577320764188 ppscbe1 = 4.33680868994202e-19
+ pscbe2 = 7.56929177375625e-08 lpscbe2 = -1.15267015861442e-13
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 4.37897997750275e-05 lalpha0 = -8.2543365127428e-11
+ alpha1 = -9.424975e-11 lalpha1 = 3.6615980750125e-16
+ beta0 = 69.7665703037275 lbeta0 = -0.000125854651189675
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.2290399268942e-09 lagidl = 1.7076707647523e-14 wagidl = 2.49248106706502e-14 pagidl = -5.25299936870593e-20
+ bgidl = 2466600645.75 lbgidl = -2349.64748473552
+ cgidl = 840.441146375 lcgidl = -0.000701012951461143
+ egidl = -1.56307736015895 legidl = 6.71638300851282e-06 wegidl = 8.470329472543e-22 pegidl = -1.61558713389263e-27
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.5769424975 lkt1 = 3.6615980750127e-9
+ kt2 = -0.019032
+ at = 472060.306850596 lat = -0.882820199830169 wat = -0.567251580053664 pat = 2.02585150855912e-6
+ ute = -1.65628748425 lute = 3.8922787537383e-7
+ ua1 = -4.7771419424e-10 lua1 = 1.94176010557143e-15 wua1 = -4.93038065763132e-32 pua1 = -1.88079096131566e-37
+ ub1 = -5.2623928494625e-18 lub1 = 4.66212205123204e-24 wub1 = 5.60547962419525e-24 pub1 = -1.81540948533207e-29
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.44 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.00636634803092+0*(0.0/sqrt(l*w*mult))} lvth0 = -4.03120386609043e-10 wvth0 = 1.58023490417281e-08 pvth0 = 2.17332616657162e-13
+ k1 = 0.55931480325 lk1 = 1.77664487477661e-8
+ k2 = 0.0221769375501519 lk2 = 1.18806290667985e-09 wk2 = -7.79000020711093e-09 pk2 = 2.40169977547548e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 167055.68835715 lvsat = -0.105461923362636 wvsat = 0.142923220740455 pvsat = -1.26486335739199e-7
+ ua = 3.42990968139568e-09 lua = -1.57329298823623e-15 wua = 1.42540012979876e-17 pua = -2.10606073322592e-23
+ ub = -3.74759715313204e-19 lub = 2.14818082619028e-24 wub = 3.0745125966889e-24 pub = -6.42024402398457e-30
+ uc = 5.181291727e-13 luc = -9.76670899893637e-19
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.025126009452831 lu0 = -2.40238443333509e-09 wu0 = 1.4364200903804e-09 pu0 = -1.50514944939576e-14
+ a0 = 1.00633244380954 la0 = -1.58104714774675e-07 wa0 = -4.97987158389925e-08 pa0 = 1.14010356013564e-13
+ keta = 0.04266318224 lketa = -1.12690999606489e-07 pketa = 5.04870979341448e-29
+ a1 = 0.0
+ a2 = 0.5
+ ags = -0.328772365208408 lags = 1.01730737639927e-06 wags = 1.38290803169269e-07 pags = -3.92434102024061e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.107717861901765+0*(0.009/sqrt(l*w*mult))} lvoff = -2.3930724238282e-08 wvoff = -1.52374500301897e-07 pvoff = 2.87225171196574e-13
+ nfactor = {0.899932471691792+0*(0.02/sqrt(l*w*mult))} lnfactor = 2.88629254704546e-07 wnfactor = -2.0381872442037e-09 pnfactor = 1.3944992028911e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.4424975e-05 lcit = -8.341055750125e-12
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.281620814262255 leta0 = -2.59791545780261e-07 weta0 = -5.5348218779072e-08 peta0 = 1.04331115657457e-13
+ etab = -0.02847850446 letab = 2.52033340545777e-8
+ dsub = 0.287980960921248 ldsub = 9.74361281825173e-09 wdsub = 3.35508411756559e-12 pdsub = -6.32431678639256e-18
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.0769779546848133 lpclm = 9.96623441931215e-07 wpclm = -1.1719704101908e-11 ppclm = 1.0371879530944e-17
+ pdiblc1 = 0.00331213796899998 lpdiblc1 = 3.50647640826125e-7
+ pdiblc2 = 0.0058837902087835 lpdiblc2 = -3.87415898724585e-9
+ pdiblcb = -0.401999 lpdiblcb = 3.33642230005e-07 wpdiblcb = -4.2351647362715e-22
+ drout = 1.52153692559705 ldrout = -9.83094497065811e-07 wdrout = 1.6940658945086e-21
+ pscbe1 = 429292893.4686 lpscbe1 = -114.883496156743
+ pscbe2 = 1.453303481712e-08 lpscbe2 = 1.90576441778914e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -6.0014119919695e-05 lalpha0 = 1.13126504477525e-10 walpha0 = -5.10787436130605e-27 palpha0 = -3.57722679260316e-32
+ alpha1 = 1.884995e-10 lalpha1 = -1.668211150025e-16
+ beta0 = -38.730102860375 lbeta0 = 7.86610352412926e-05 wbeta0 = 1.35525271560688e-20 pbeta0 = 3.87740912134232e-26
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 6.82979960568214e-09 lagidl = 6.51930365680616e-15 wagidl = 1.63242721513103e-14 pagidl = -3.63180215807962e-20
+ bgidl = 915927218.5 lbgidl = 573.364172263592
+ cgidl = 1295.31598933932 lcgidl = -0.00155844975607467 wcgidl = -0.00370401286624304 pcgidl = 6.9820457328038e-9
+ egidl = 3.0805973382958 legidl = -2.03692057970089e-6
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.526325275 lkt1 = -9.17516132513746e-8
+ kt2 = -0.019032
+ at = -19538.7317183299 lat = 0.0438415298770634 wat = 0.956585116415867 pat = -8.46573045102461e-7
+ ute = -1.440065055 lute = -1.83503226502754e-8
+ ua1 = 5.524e-10
+ ub1 = -2.07953361254055e-18 lub1 = -1.33755169606968e-24 wub1 = -7.58779378911078e-24 pub1 = 6.71515956439409e-30
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.81e-6
+ sbref = 2.81e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.45 pmos
* DC IV MOS Parameters
+ lmin = 8.0e-07 lmax = 1e-06 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.28260034036115+0*(0.0/sqrt(l*w*mult))} lvth0 = 2.44062581655683e-07 wvth0 = 1.15658808273674e-06 pvth0 = -7.92257053734256e-13
+ k1 = 0.5898704235 lk1 = -9.27512239538251e-9
+ k2 = -0.0119116721231175 lk2 = 3.13563120244748e-08 wk2 = 8.56144326073133e-08 pk2 = -5.86454582638466e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 7759.59541750001 lvsat = 0.0355143224084896
+ ua = -7.21237315312302e-10 lua = 2.10045134811535e-15 wua = -4.22294372677093e-17 pua = 2.89269533811939e-23
+ ub = 9.86620178993335e-18 lub = -6.91501890114539e-24 wub = -1.84965787423894e-23 pub = 1.2670063955643e-29
+ uc = 5.8546574915e-12 luc = -5.69947177939004e-18 wuc = 3.08148791101958e-33
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0344640438218651 lu0 = -1.06664981597585e-08 wu0 = -6.89013494803565e-08 pu0 = 4.71970798872969e-14
+ a0 = 0.773471669422749 la0 = 4.79759062537641e-08 wa0 = 3.49693707448171e-07 pa0 = -2.39538441133458e-13
+ keta = -0.15139736295 lketa = 5.90516125839353e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 1.16190941325825 lags = -3.01938544134836e-07 wags = -1.35023716336637e-06 pags = 9.24905705720148e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.346891229018449+0*(0.009/sqrt(l*w*mult))} lvoff = 1.87736509793147e-07 wvoff = 7.61872501509483e-07 pvoff = -5.21878854171489e-13
+ nfactor = {-0.597322326302884+0*(0.02/sqrt(l*w*mult))} lnfactor = 1.61369226465584e-06 wnfactor = 6.96347708685455e-06 pnfactor = -4.76994698710994e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -1.2124875e-05 lcit = 1.5155428750625e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -0.055229775771966 leta0 = 3.83195421470748e-08 weta0 = 2.7674109389536e-07 peta0 = -1.89566265612852e-13
+ etab = 0.001821812702 letab = -1.61229513220649e-9
+ dsub = 0.381762965481509 ldsub = -7.32529923075563e-08 wdsub = -1.67754205878279e-11 pdsub = 1.14910792264315e-17
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.99395583862875 lpclm = -6.9989240046975e-7
+ pdiblc1 = 0.20282696902275 lpdiblc1 = 1.74078012917711e-7
+ pdiblc2 = -0.0324173066339675 lpdiblc2 = 3.00221202131046e-08 wpdiblc2 = -1.98523347012727e-23 ppdiblc2 = -6.31088724176809e-30
+ pdiblcb = -0.025
+ drout = 0.3384020931485 ldrout = 6.39739139769935e-8
+ pscbe1 = -44797159.5074992 lpscbe1 = 304.68383027684
+ pscbe2 = 1.815406017615e-08 lpscbe2 = -3.18553169343688e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.00024102438742525 lalpha0 = -1.53291069330214e-10
+ alpha1 = 0.0
+ beta0 = 66.614022720125 lbeta0 = -1.4567989176822e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 5.60057844418412e-09 lagidl = 7.60715823862608e-15 wagidl = -1.09355611741237e-13 pagidl = 7.49080472646886e-20
+ bgidl = 729818587.499998 lbgidl = 738.069380155437
+ cgidl = -3841.4949104466 lcgidl = 0.00298760220618137 wcgidl = 0.0185200643312152 pcgidl = -1.26861514665608e-8
+ egidl = 1.79942371219525 legidl = -9.03088326470036e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.5940377625 lkt1 = -3.18264003763125e-8
+ kt2 = -0.019032
+ at = 47124.875 lat = -0.015155428750625
+ ute = -1.395725475 lute = -5.75906292523759e-8
+ ua1 = 5.524e-10
+ ub1 = -3.5909e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.41e-6
+ sbref = 2.41e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.46 pmos
* DC IV MOS Parameters
+ lmin = 6e-07 lmax = 8.0e-07 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.643958083601703+0*(0.0/sqrt(l*w*mult))} lvth0 = -1.93404171013252e-07 wvth0 = -1.0584980245721e-06 pvth0 = 7.25065854341761e-13
+ k1 = 0.619488790519179 lk1 = -2.95635557116849e-08 wk1 = -1.30360522540111e-07 pk1 = 8.92963061373642e-14
+ k2 = 0.0166312130745965 lk2 = 1.18045783784668e-08 wk2 = 2.33508975494986e-09 pk2 = -1.59952480669181e-15
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 110685.785476972 lvsat = -0.0349896031512983 wvsat = -0.252866317967508 pvsat = 1.73212163476153e-7
+ ua = -8.12643544951376e-09 lua = 7.17297504405268e-15 wua = 3.16296010253265e-14 pua = -2.16661185543435e-20
+ ub = 5.98459175947591e-18 lub = -4.2561354383322e-24 wub = -1.79812097270695e-23 pub = 1.2317038756994e-29
+ uc = 1.00812943608082e-11 luc = -8.59469690168182e-18 wuc = -3.78983228575002e-17 puc = 2.59601616657733e-23
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = -0.017623841894412 lu0 = 2.50134431164627e-08 wu0 = 1.21163578481639e-07 pu0 = -8.29964454420304e-14
+ a0 = 1.07196548775526 la0 = -1.56490866834911e-07 wa0 = -6.90046602387919e-07 pa0 = 4.72678472402711e-13
+ keta = 0.209042887964679 lketa = -1.87848157091365e-07 wketa = -9.90666425170827e-07 pketa = 6.78601547909891e-13
+ a1 = 0.0
+ a2 = 0.5
+ ags = -2.49831880532906 lags = 2.20529948445638e-06 wags = 9.72426983935314e-06 pags = -6.6610762186077e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {0.128341298540492+0*(0.009/sqrt(l*w*mult))} lvoff = -1.37795395422089e-07 wvoff = -6.07608906250242e-07 pvoff = 4.16209062736885e-13
+ nfactor = {2.2089329937628+0*(0.02/sqrt(l*w*mult))} lnfactor = -3.08578598312547e-07 wnfactor = -2.57245990248053e-06 pnfactor = 1.76212217089965e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -0.141012283472997 leta0 = 9.70801310097426e-08 weta0 = 4.31514841851966e-07 peta0 = -2.95585509094387e-13
+ etab = -0.001821812702 letab = 8.8357005140649e-10
+ dsub = 0.07042821565198 ldsub = 1.40009754651922e-07 wdsub = 6.17398834400736e-07 pdsub = -4.22915114570332e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.822013671729616 lpclm = 1.22903263427818e-06 wpclm = 5.41940317036867e-06 ppclm = -3.71226407468668e-12
+ pdiblc1 = -0.21387973730657 lpdiblc1 = 4.59520023219763e-07 wpdiblc1 = 2.02625390967083e-06 ppdiblc1 = -1.38797379685497e-12
+ pdiblc2 = 0.0480005979750318 lpdiblc2 = -2.50637423545369e-08 wpdiblc2 = -1.10518591945176e-07 ppdiblc2 = 7.57046828894859e-14
+ pdiblcb = -0.025
+ drout = -2.36559029483992 ldrout = 1.91619517978712e-06 wdrout = 8.44946417683997e-06 pdrout = -5.78784071381449e-12
+ pscbe1 = 477038380.203968 lpscbe1 = -52.7709052478169 wpscbe1 = -232.693348868763 ppscbe1 = 0.000159393780508358
+ pscbe2 = 6.43200760613525e-09 lpscbe2 = 4.84401570676037e-15 wpscbe2 = 2.13596911306649e-14 ppscbe2 = -1.46312816260498e-20
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -0.000314774225878372 lalpha0 = 2.274282017897e-10 walpha0 = 1.00284483756957e-09 palpha0 = -6.86943699510965e-16
+ alpha1 = 0.0
+ beta0 = 0.208758917117564 lbeta0 = 3.09192845019191e-05 wbeta0 = 0.000136338609724251 pbeta0 = -9.33912659680635e-11
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 6.03488474047472e-08 lagidl = -2.98951322580148e-14 wagidl = -9.51116991604709e-14 pagidl = 6.51510383664268e-20
+ bgidl = 2416636379.54439 lbgidl = -417.392373306011 wbgidl = -1840.49200370452 pbgidl = 0.00126072782007758
+ cgidl = 2285.31019048825 lcgidl = -0.0012092286539335 wcgidl = -0.00533209471602709 pcgidl = 3.65245822000498e-9
+ egidl = -1.25886005847704 legidl = 1.19182076502163e-06 wegidl = 5.25533461595651e-06 pegidl = -3.59987793525713e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.792780090510974 lkt1 = 1.04311100599566e-07 wkt1 = 4.96436404595627e-07 pkt1 = -3.40056454965981e-13
+ kt2 = -0.019032
+ at = 41974.825 lat = -0.011627670250875
+ ute = -1.71698023306775 lute = 1.62467273750243e-07 wute = 5.51596005106252e-07 pute = -3.77840505517757e-13
+ ua1 = 5.53369990000001e-10 lua1 = -6.64438300049995e-19
+ ub1 = -4.2982652075e-18 lub1 = 4.84541630311463e-25
+ uc1 = -2.733805074e-10 luc1 = 1.12462826666463e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.02e-6
+ sbref = 2.01e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.47 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 6e-07 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.02/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.10393502170036+0*(0.0/sqrt(l*w*mult))} lvth0 = 2.96823440799076e-08 wvth0 = 1.19828503443329e-06 pvth0 = -3.69462645360557e-13
+ k1 = 0.348851753494348 lk1 = 1.01694054060173e-07 wk1 = 7.75356844249433e-07 pk1 = -3.49972088168731e-13
+ k2 = 0.0779599527519153 lk2 = -1.79395537213344e-08 wk2 = -1.8676309585803e-07 pk2 = 9.01121497246755e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 164525.831571966 lvsat = -0.0611017563071399 wvsat = -0.742041704747214 pvsat = 4.10459780187377e-7
+ ua = 2.0059489251961e-08 lua = -6.49705750653907e-15 wua = -5.64206325861463e-14 pua = 2.10378044960527e-20
+ ub = -1.50400468993476e-17 lub = 5.94070918800392e-24 wub = 3.98153280833134e-23 pub = -1.57139930983527e-29
+ uc = -1.51198930834481e-10 luc = 6.96254059169073e-17 wuc = 8.39206164184256e-16 puc = -3.99431129027043e-22
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0662423922121323 lu0 = -1.56612610940407e-08 wu0 = -1.71612169811411e-07 pu0 = 5.89983286013574e-14
+ a0 = 1.29663151009379 la0 = -2.65452764338988e-07 wa0 = -2.32510940376347e-06 pa0 = 1.26567575575585e-12
+ keta = -0.138825918894737 lketa = -1.91335251085827e-08 wketa = -2.00482405011294e-07 pketa = 2.95366249052618e-13
+ a1 = 0.0
+ a2 = 0.5
+ ags = -1.03938558546288 lags = 1.49772416748738e-06 wags = 1.14938282804182e-05 pags = -7.51930321473207e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.170704255016395+0*(0.009/sqrt(l*w*mult))} lvoff = 7.24020282523301e-09 wvoff = 8.49086989259772e-07 pvoff = -2.90281163105995e-13
+ nfactor = {6.13865940944519+0*(0.02/sqrt(l*w*mult))} lnfactor = -2.21447626128643e-06 wnfactor = -1.29563654511268e-05 pnfactor = 6.79826444246534e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 5.832155018925e-05 lcit = -2.34357102340353e-11 wcit = -1.45954565844927e-10 pcit = 7.07872346619603e-17
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.733271128413976 leta0 = -3.2694295233838e-07 weta0 = -3.88350104203835e-06 peta0 = 1.797175619513e-12
+ etab = 0.0110128759253299 letab = -5.34118975940538e-09 wetab = 1.4242246535148e-07 petab = -6.90741835831408e-14
+ dsub = 0.638774274315756 ldsub = -1.35635242069716e-07 wdsub = -1.31247322919848e-06 pdsub = 5.13063186914971e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.380902234560436 lpclm = 6.45624434307035e-07 wpclm = 6.04819530934705e-06 ppclm = -4.01722511813051e-12
+ pdiblc1 = 0.86364312659068 lpdiblc1 = -6.3073178156083e-08 wpdiblc1 = 1.88374402251968e-06 ppdiblc1 = -1.3188572141361e-12
+ pdiblc2 = -0.0725936641882034 lpdiblc2 = 3.34238718233214e-08 wpdiblc2 = 3.41908272443753e-07 ppdiblc2 = -1.43720084204823e-13
+ pdiblcb = -1.18787200757 lpdiblcb = 5.63987109311411e-07 wpdiblcb = 5.83818263379707e-06 ppdiblcb = -2.83148938647841e-12
+ drout = 6.51925799190087 ldrout = -2.39291181504073e-06 wdrout = -2.49945885059457e-05 pdrout = 1.04323576170731e-11
+ pscbe1 = 858383169.460168 lpscbe1 = -237.721221313128 wpscbe1 = -1016.4511853715 ppscbe1 = 0.000539512412423004
+ pscbe2 = 2.44556428481255e-08 lpscbe2 = -3.89735726742868e-15 wpscbe2 = -4.51688501671656e-14 ppscbe2 = 1.76347282606915e-20
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.000321626784423965 lalpha0 = -8.12231062018815e-11 walpha0 = -7.18915544690304e-10 palpha0 = 1.48101477083161e-16
+ alpha1 = 5.81436003784999e-10 lalpha1 = -2.81993554655706e-16 walpha1 = -2.91909131689854e-15 palpha1 = 1.41574469323921e-21
+ beta0 = -160.728224917988 lbeta0 = 0.000108972916977026 wbeta0 = 0.00111488478557166 pbeta0 = -5.67981268523178e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -2.39229444728862e-08 lagidl = 1.0976265443678e-14 wagidl = 5.40185974744559e-14 pagidl = -7.17640985002951e-21
+ bgidl = -1516050963.18562 lbgidl = 1489.94132448133 wbgidl = 16866.5194858397 pbgidl = -0.00781207921729394
+ cgidl = -406.499855831804 lcgidl = 9.62857594814959e-05 wcgidl = -9.0326797663411e-05 pcgidl = 1.11022698843818e-9
+ egidl = 10.9245997905903 legidl = -4.7170963444768e-06 wegidl = -4.92082311709207e-05 pegidl = 2.28146791535494e-11
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.590350128205151 lkt1 = 6.13358103105179e-09 wkt1 = -8.17727330177337e-07 pkt1 = 2.97306385580233e-13
+ kt2 = -0.019032
+ at = 18000.0
+ ute = -0.837488160079502 lute = -2.64081984188693e-07 wute = -4.02228332711104e-06 pute = 1.84046810121097e-12
+ ua1 = 5.52e-10
+ ub1 = -4.85919974e-18 lub1 = 7.565920739013e-25
+ uc1 = -4.1496e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 1.81e-6
+ sbref = 1.81e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.48 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 1.5e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.983061556614667+0*(0.0/sqrt(l*w*mult))} wvth0 = 8.06063706428084e-8
+ k1 = 0.609218744346667 wk1 = -4.23132161766861e-8
+ k2 = 0.0192169592623827 wk2 = 7.67819845940281e-9
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 219918.3666 wvsat = -0.0601631474581675
+ ua = 2.7300353730846e-09 wua = -7.75338279860369e-17
+ ub = -1.26132060933333e-19 wub = -3.09235516197197e-26
+ uc = -5.65199559666667e-11 wuc = 4.99828693259331e-17
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0206626855638533 wu0 = -1.2835723312411e-9
+ a0 = 0.829738468194666 wa0 = 1.97108555066764e-7
+ keta = -0.00620795355146667 wketa = -5.18903319654465e-9
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.125356374758693 wags = 2.77236069920134e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0873158714868107+0*(0.009/sqrt(l*w*mult))} wvoff = -1.77869941995912e-8
+ nfactor = {1.90324784953333+0*(0.02/sqrt(l*w*mult))} wnfactor = -3.8287030990554e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.50682866666667e-05 wcit = -1.53086889206533e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.0800000000000101
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.68498419736076 wpclm = 2.32129014953691e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00461412075788147 wpdiblc2 = -5.05427907466816e-9
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 450686940.044587 wpscbe1 = -353.318661752133
+ pscbe2 = 1.501696871758e-08 wpscbe2 = -4.83601483003367e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 8.16002977865213e-05 walpha0 = -9.34330220261647e-11
+ alpha1 = 0.0
+ beta0 = 39.0737200539413 wbeta0 = -2.43956817249307e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.98179452333333e-08 wagidl = -1.52321454760501e-14
+ bgidl = 1758467825.33333 wbgidl = 52.0495423302227
+ cgidl = 1539.26570133333 wcgidl = -0.00162884450115751
+ egidl = 0.49239983118232 wegidl = 6.07445163520939e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.555726853333333 wkt1 = -6.12347556826136e-8
+ kt2 = -0.019032
+ at = 557494.475853333 wat = -0.328310142592332
+ ute = -1.51582685333333 wute = -6.12347556826132e-8
+ ua1 = 2.2096e-11
+ ub1 = -3.5705585484e-18 wub1 = -2.78311964577476e-25
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.49 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 1.5e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.983061556614667+0*(0.0/sqrt(l*w*mult))} wvth0 = 8.06063706428079e-8
+ k1 = 0.609218744346667 wk1 = -4.23132161766861e-8
+ k2 = 0.0192169592623827 wk2 = 7.67819845940284e-9
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 219918.3666 wvsat = -0.0601631474581675
+ ua = 2.7300353730846e-09 wua = -7.75338279860369e-17
+ ub = -1.26132060933333e-19 wub = -3.09235516197198e-26
+ uc = -5.65199559666667e-11 wuc = 4.99828693259332e-17
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0206626855638533 wu0 = -1.28357233124111e-9
+ a0 = 0.829738468194666 wa0 = 1.97108555066764e-7
+ keta = -0.00620795355146667 wketa = -5.18903319654465e-9
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.125356374758693 wags = 2.77236069920135e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0873158714868106+0*(0.009/sqrt(l*w*mult))} wvoff = -1.77869941995912e-8
+ nfactor = {1.90324784953333+0*(0.02/sqrt(l*w*mult))} wnfactor = -3.82870309905539e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.50682866666667e-05 wcit = -1.53086889206533e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.0800000000000101
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.68498419736076 wpclm = 2.32129014953691e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00461412075788147 wpdiblc2 = -5.05427907466816e-9
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 450686940.044587 wpscbe1 = -353.318661752133
+ pscbe2 = 1.501696871758e-08 wpscbe2 = -4.83601483003367e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 8.16002977865213e-05 walpha0 = -9.34330220261647e-11
+ alpha1 = 0.0
+ beta0 = 39.0737200539413 wbeta0 = -2.43956817249304e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.98179452333333e-08 wagidl = -1.52321454760501e-14
+ bgidl = 1758467825.33333 wbgidl = 52.0495423302218
+ cgidl = 1539.26570133333 wcgidl = -0.00162884450115751
+ egidl = 0.49239983118232 wegidl = 6.07445163520939e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.555726853333333 wkt1 = -6.12347556826136e-8
+ kt2 = -0.019032
+ at = 557494.475853333 wat = -0.328310142592331
+ ute = -1.51582685333333 wute = -6.12347556826123e-8
+ ua1 = 2.2096e-11
+ ub1 = -3.5705585484e-18 wub1 = -2.78311964577476e-25
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.50 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 1.5e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.994379552280467+0*(0.0/sqrt(l*w*mult))} lvth0 = 8.92423392348648e-08 wvth0 = 9.78152246007195e-08 pvth0 = -1.35691727413864e-13
+ k1 = 0.627113968183211 lk1 = -1.41103750475031e-07 wk1 = -6.95226534870179e-08 pk1 = 2.14546277144779e-13
+ k2 = 0.0149942731656086 lk2 = 3.3295858759633e-08 wk2 = 1.40987335519425e-08 pk2 = -5.06258871019994e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 366776.547789739 lvsat = -1.15797602439018 wvsat = -0.283458955942628 pvsat = 1.76068633342093e-6
+ ua = 2.22053586114902e-09 lua = 4.01740110411452e-15 wua = 6.97153046918854e-16 pua = -6.10840213519067e-21
+ ub = 3.74073671136017e-19 lub = -3.94411969633817e-24 wub = -7.91479364350918e-25 pub = 5.99697878060644e-30
+ uc = -7.97407201864798e-11 luc = 1.83095609769405e-16 wuc = 8.52897162314599e-17 puc = -2.78394311315844e-22
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0192264325005918 lu0 = 1.13248482225519e-08 wu0 = 9.00230343905172e-10 pu0 = -1.7219273174515e-14
+ a0 = 0.867476366046469 la0 = -2.97563135871976e-07 wa0 = 1.39728609713667e-07 pa0 = 4.52440582209438e-13
+ keta = -0.000266152509083593 lketa = -4.68510715101853e-08 wketa = -1.42234584962735e-08 pketa = 7.12363983162356e-14
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.0843231154420394 lags = 3.2354704454552e-07 wags = 9.01141033173553e-08 pags = -4.91948751572839e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0904613433391115+0*(0.009/sqrt(l*w*mult))} lvoff = 2.48020298280327e-08 wvoff = -1.30043482847736e-08 pvoff = -3.77111391251059e-14
+ nfactor = {1.89448603502101+0*(0.02/sqrt(l*w*mult))} lnfactor = 6.90868636205636e-08 wnfactor = -3.69548093604962e-07 pnfactor = -1.05045608918975e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.50682866666667e-05 wcit = -1.53086889206533e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.0800000000000101
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -2.14953678715502 lpclm = 1.15479898477648e-05 wpclm = 4.54812185858283e-06 ppclm = -1.75585568916685e-11
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0078426688888229 lpdiblc2 = -2.54570858697325e-08 wpdiblc2 = -9.96324130809077e-09 ppdiblc2 = 3.87071426657261e-14
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 907773651.118053 lpscbe1 = -3604.12643138073 wpscbe1 = -1048.31260672538 ppscbe1 = 0.00548002378114435
+ pscbe2 = -4.5655002089364e-08 lpscbe2 = 4.78398186452899e-13 wpscbe2 = 9.22025220560667e-14 ppscbe2 = -7.27397744927023e-19
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.000136604348573555 lalpha0 = -4.33706665435503e-10 walpha0 = -1.77065911191138e-10 palpha0 = 6.59444912901367e-16
+ alpha1 = 0.0
+ beta0 = 40.8232216763534 lbeta0 = -1.37948115452114e-05 wbeta0 = -5.09966089634796e-06 pbeta0 = 2.09748178271322e-11
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 3.03301668859481e-08 lagidl = -8.28888151697594e-14 wagidl = -3.12158313277477e-14 pagidl = 1.26031283022207e-19
+ bgidl = 1590076702.6747 lbgidl = 1327.76316020768 wbgidl = 308.085886856952 pbgidl = -0.00201884529641153
+ cgidl = 2204.22483842897 lcgidl = -0.00524319947120338 wcgidl = -0.00263990555968351 pcgidl = 7.97221139117215e-9
+ egidl = 1.52462112158086 legidl = -8.13905971368604e-06 wegidl = -9.62032857431976e-07 pegidl = 1.23753263478236e-11
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.555726853333333 wkt1 = -6.12347556826132e-8
+ kt2 = -0.019032
+ at = 986080.197333148 lat = -3.37939627093973 wat = -0.979968731902289 pat = 5.13832471841607e-6
+ ute = -1.47671160997477 lute = -3.08423498306083e-07 wute = -1.20708935595907e-07 pute = 4.6895361124542e-13
+ ua1 = 2.2096e-11
+ ub1 = -3.39277976733532e-18 lub1 = -1.40178479980115e-24 wub1 = -5.48622112283399e-25 pub1 = 2.13139416311044e-30
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.51 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 1.5e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.943092723348517+0*(0.0/sqrt(l*w*mult))} lvth0 = -1.1000673473162e-07 wvth0 = 1.3199278030269e-08 pvth0 = 1.93040801932606e-13
+ k1 = 0.623664836230371 lk1 = -1.27703890083908e-07 wk1 = -6.42782966405716e-08 pk1 = 1.94171977018121e-13
+ k2 = 0.0205853441726288 lk2 = 1.15745758527145e-08 wk2 = 8.56257761184345e-09 pk2 = -2.91179489554946e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 47266.9403114863 lvsat = 0.0833172031147901 wvsat = 0.202350929093549 pvsat = -1.26682640895195e-7
+ ua = 3.9537492448964e-09 lua = -2.71612422567715e-15 wua = -1.93757321701042e-15 pua = 4.12749622654324e-21
+ ub = -2.56589743296638e-18 lub = 7.47765334324412e-24 wub = 3.58451088374003e-24 pub = -1.10037214532757e-29
+ uc = -9.82948057585349e-11 luc = 2.55178139446412e-16 wuc = 1.32033201196519e-16 puc = -4.59992516687675e-22
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0209471143013298 lu0 = 4.64000803009386e-09 wu0 = -1.94977339336402e-09 pu0 = -6.14702290524283e-15
+ a0 = 0.602467981646854 la0 = 7.31993112478605e-07 wa0 = 6.82115211905555e-07 pa0 = -1.65472865537303e-12
+ keta = -0.000642376628333031 lketa = -4.53894426880219e-08 wketa = -1.36514149900924e-08 pketa = 6.90140121549396e-14
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.0949743178810095 lags = 2.82167176326133e-07 wags = 9.10322890914152e-08 pags = -4.95515898714133e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0293866559210917+0*(0.009/sqrt(l*w*mult))} lvoff = -2.12472825417537e-07 wvoff = -1.05867555458249e-07 pvoff = 3.23061956427809e-13
+ nfactor = {2.74616461449315+0*(0.02/sqrt(l*w*mult))} lnfactor = -3.23968015923577e-06 wnfactor = -1.53844766748676e-06 pnfactor = 4.43612339111395e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.50682866666667e-05 wcit = -1.53086889206533e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -0.0410839147609786 leta0 = 4.70410403426867e-07 weta0 = 1.84106397219277e-07 peta0 = -7.15252432664904e-13
+ etab = -0.174177715502511 letab = 4.04729903838677e-07 wetab = 1.58400757933551e-07 petab = -6.15386152568055e-13
+ dsub = 1.06644580962335 ldsub = -1.96753943815767e-06 wdsub = -7.70043763290971e-07 pdsub = 2.99161617016661e-12
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.25313312052394 lpclm = -1.6713657302184e-06 wpclm = -6.25590098664317e-07 ppclm = 2.54128819367686e-12
+ pdiblc1 = 0.770840036942151 lpdiblc1 = -1.47956163932007e-06 wpdiblc1 = -5.79061944410023e-07 ppdiblc1 = 2.24965275872322e-12
+ pdiblc2 = -0.00352778852618155 lpdiblc2 = 1.87170843352727e-08 wpdiblc2 = 7.32538000501969e-09 ppdiblc2 = -2.84590646926015e-14
+ pdiblcb = 0.354573400504667 lpdiblcb = -1.47464076309363e-06 wpdiblcb = -5.77136041439739e-07 ppdiblcb = 2.24217063531318e-12
+ drout = -0.275061481110266 ldrout = 3.24420967880598e-06 wdrout = 1.26969929116743e-06 pdrout = -4.93277539768899e-12
+ pscbe1 = -529216733.400988 lpscbe1 = 1978.57402752383 wpscbe1 = 1136.61115507043 ppscbe1 = -0.00300839410881359
+ pscbe2 = 1.37229778517494e-07 lpscbe2 = -2.32108271780842e-13 wpscbe2 = -1.85871226469733e-13 ppscbe2 = 3.52917377726965e-19
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 6.77515925394678e-05 lalpha0 = -1.66214052506856e-10 walpha0 = -7.23762595798933e-11 palpha0 = 2.5272613983994e-16
+ alpha1 = -1.89786700252333e-10 lalpha1 = 7.37320381546814e-16 walpha1 = 2.88568020719869e-16 palpha1 = -1.12108531765659e-21
+ beta0 = 102.504981821987 lbeta0 = -0.000253428141302197 wbeta0 = -9.88859136531419e-05 pbeta0 = 3.85333940856013e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.89023327679214e-08 lagidl = -3.84917367603962e-14 wagidl = -2.84571229295728e-14 pagidl = 1.15313714688839e-19
+ bgidl = 2966369569.71833 lbgidl = -4019.12774679247 wbgidl = -1509.5450380814 pbgidl = 0.00504264175881934
+ cgidl = 1917.29932148017 lcgidl = -0.0041284952724849 wcgidl = -0.00325263504189072 pcgidl = 1.03526623658998e-8
+ egidl = -4.05159033100872 legidl = 1.35244938985672e-05 wegidl = 7.51651858927015e-06 pegidl = -2.05638036298569e-11
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.551892503320716 lkt1 = -1.48964306272656e-08 wkt1 = -7.56631567186068e-08 pkt1 = 5.60542658828294e-14
+ kt2 = -0.019032
+ at = 178329.6922915 lat = -0.241289597605455 wat = 0.319957628993481 pat = 8.8117305967808e-8
+ ute = -1.61807270414907 lute = 2.40763645755603e-07 wute = -1.15427208287947e-07 pute = 4.48434127062635e-13
+ ua1 = -4.7771419424e-10 lua1 = 1.94176010557143e-15 pua1 = -9.4039548065783e-38
+ ub1 = -3.53182136228081e-18 lub1 = -8.61608898645871e-25 wub1 = 3.7831267516375e-25 pub1 = -1.46974285144779e-30
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.52 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 1.5e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.06553521189804+0*(0.0/sqrt(l*w*mult))} lvth0 = 1.20796743971791e-07 wvth0 = 1.94521073988289e-07 pvth0 = -1.48749876839283e-13
+ k1 = 0.536938118179587 lk1 = 3.57755398082304e-08 wk1 = 6.75884639815932e-08 pk1 = -5.43962074208567e-14
+ k2 = 0.0175957238521783 lk2 = 1.72099952086623e-08 wk2 = 6.04749163062668e-09 pk2 = -2.43770244563309e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 221949.50887766 lvsat = -0.245958565219605 wvsat = -0.0228827956282576 pvsat = 2.97881804036788e-7
+ ua = 4.20120455293167e-09 lua = -3.18257624404709e-15 wua = -2.31543136004826e-15 pua = 4.83975693687886e-21
+ ub = 1.35805036428499e-18 lub = 8.10313651642732e-26 wub = -2.15941598939634e-24 pub = -1.76448017047973e-31
+ uc = 6.96236467717724e-11 luc = -6.1347303980955e-17 wuc = -2.08732248430752e-16 puc = 1.82348652032483e-22
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0311859048221171 lu0 = -1.46600609076376e-08 wu0 = -1.68674090340131e-08 pu0 = 2.19726456892025e-14
+ a0 = 1.13080406676251 la0 = -2.63917766283977e-07 wa0 = -4.25763510365708e-07 pa0 = 4.33617196714689e-13
+ keta = 0.0956611228877124 lketa = -2.2692105775827e-07 wketa = -1.60079537755246e-07 pketa = 3.45030291426641e-13
+ a1 = 0.0
+ a2 = 0.5
+ ags = -0.740635177276849 lags = 1.85728689665122e-06 wags = 1.38231666094263e-06 pags = -2.92958048323181e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.218123493168684+0*(0.009/sqrt(l*w*mult))} lvoff = 1.43295169109988e-07 wvoff = 1.81104163260994e-07 pvoff = -2.17878298499369e-13
+ nfactor = {0.190001023648461+0*(0.02/sqrt(l*w*mult))} lnfactor = 1.5786754286885e-06 wnfactor = 2.1422998125304e-06 pnfactor = -2.50206720498101e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 2.39786700252333e-05 lcit = -1.67960280789814e-11 wcit = -2.88568020719869e-11 pcit = 2.55381255496981e-17
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.449096418672437 leta0 = -4.53577074193454e-07 weta0 = -5.61205937241563e-07 peta0 = 6.89657591232108e-13
+ etab = 0.0136100639850883 letab = 5.07508784434501e-08 wetab = -1.27127931748431e-07 petab = -7.71660001609677e-14
+ dsub = 0.0122491038755299 ldsub = 1.96160811934424e-08 wdsub = 8.32847569044711e-07 pdsub = -2.98259768294925e-14
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.698190111128697 lpclm = 2.00686880483065e-06 wpclm = 2.34137257073268e-06 ppclm = -3.05142160332315e-12
+ pdiblc1 = -0.388656849089711 lpdiblc1 = 7.06084193365559e-07 wpdiblc1 = 1.18393683784502e-06 ppdiblc1 = -1.07359113083363e-12
+ pdiblc2 = 0.0105403193417118 lpdiblc2 = -7.80122865516685e-09 wpdiblc2 = -1.40649810546019e-08 ppdiblc2 = 1.186165895298e-14
+ pdiblcb = -0.784146801009333 lpdiblcb = 6.71841123159255e-07 wpdiblcb = 1.15427208287948e-06 ppdiblcb = -1.02152502198792e-12
+ drout = 2.49620588149929 ldrout = -1.97961544337622e-06 wdrout = -2.94397393593733e-06 pdrout = 3.00997756703733e-12
+ pscbe1 = 643152435.768598 lpscbe1 = -231.335994514999 wpscbe1 = -645.959753483553 ppscbe1 = 0.000351743140956132
+ pscbe2 = 1.4074731768937e-08 lpscbe2 = 3.83755649548618e-17 wpscbe2 = 1.38429794079404e-15 ppscbe2 = -5.83495092559441e-23
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -0.000141273931582555 lalpha0 = 2.27798015335535e-10 walpha0 = 2.45444123490304e-10 palpha0 = -3.46363693145467e-16
+ alpha1 = 3.79573400504667e-10 lalpha1 = -3.35920561579627e-16 walpha1 = -5.77136041439739e-16 palpha1 = 5.10762510993961e-22
+ beta0 = -115.970139737178 lbeta0 = 0.000158396370461221 wbeta0 = 0.000233302450025866 pbeta0 = -2.40839463737099e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -2.63465954397819e-09 lagidl = 2.10538606257297e-15 wagidl = 4.49115385104312e-14 pagidl = -2.29858452822613e-20
+ bgidl = 205822555.542801 lbgidl = 1184.48957219333 wbgidl = 2144.86119299694 pbgidl = -0.00184589571473217
+ cgidl = -1637.18713306077 lcgidl = 0.0025716939218925 wcgidl = 0.00515357175992272 pcgidl = -5.49299542448456e-9
+ egidl = 5.29917927914914 legidl = -4.10166006273228e-06 wegidl = -6.70119569220034e-06 pegidl = 6.23651670214356e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.4707517397729 lkt1 = -1.67846364211083e-07 wkt1 = -1.67859085123963e-07 pkt1 = 2.29843129947283e-13
+ kt2 = -0.019032
+ at = 50369.497281294 lat = -8.52698121922568e-05 wat = 0.745428289437709 pat = -7.1389276161626e-7
+ ute = -1.45369889818193 lute = -6.9080156623414e-08 wute = 4.11808324572238e-08 pute = 1.53228753298187e-13
+ ua1 = 5.524e-10
+ ub1 = -4.34114596193838e-18 lub1 = 6.63963925085658e-25 wub1 = -7.56625350327497e-25 pub1 = 6.69609651913085e-31
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.81e-6
+ sbref = 2.81e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.53 pmos
* DC IV MOS Parameters
+ lmin = 8.0e-07 lmax = 1e-06 wmin = 1.5e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.731640799145659+0*(0.0/sqrt(l*w*mult))} lvth0 = -1.74698141842004e-07 wvth0 = -5.07577498071057e-07 pvth0 = 4.72603848940378e-13
+ k1 = 0.583086809928764 lk1 = -5.0658216463329e-09 wk1 = 2.04898098213287e-08 pk1 = -1.27141339822935e-14
+ k2 = 0.0480867670710105 lk2 = -9.77442558478821e-09 wk2 = -9.56100130004014e-08 pk2 = 6.55893588546059e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -464784.737438231 lvsat = 0.361797809098727 wvsat = 1.42731354177007 pvsat = -9.85534703579049e-7
+ ua = -8.73528875898114e-09 lua = 8.26615565452918e-15 wua = 2.41641007516138e-14 pua = -1.85944965842815e-20
+ ub = 1.03281570561032e-17 lub = -7.8574682065614e-24 wub = -1.98919081564817e-23 pub = 1.55167188883618e-29
+ uc = 1.17910463110508e-11 luc = -1.01657417362187e-17 wuc = -1.79307793200096e-17 puc = 1.34903058768216e-23
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = -0.0111693967085531 lu0 = 2.28241691704978e-08 wu0 = 6.89338187736042e-08 pu0 = -5.39610119143998e-14
+ a0 = 0.63028205795396 la0 = 1.79041708901544e-07 wa0 = 7.82195924235083e-07 pa0 = -6.35420863109839e-13
+ keta = -0.486043777953836 lketa = 2.87884870961996e-07 wketa = 1.01079481146928e-06 pketa = -6.91187653265315e-13
+ a1 = 0.0
+ a2 = 0.5
+ ags = 3.5900678278454 lags = -1.97536360936694e-06 wags = -8.68445566040903e-06 pags = 5.9794626873028e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0367771365927949+0*(0.009/sqrt(l*w*mult))} lvoff = -1.71954497278907e-08 wvoff = -1.7482277306491e-07 pvoff = 9.71152605143735e-14
+ nfactor = {2.62819232721602+0*(0.02/sqrt(l*w*mult))} lnfactor = -5.79111684012264e-07 wnfactor = -2.77914476689413e-06 pnfactor = 1.8533866405868e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -1.2124875e-05 lcit = 1.5155428750625e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -0.261860525743615 leta0 = 1.7561626683003e-07 weta0 = 9.00866381354225e-07 peta0 = -6.04269100363572e-13
+ etab = 0.303432007034191 letab = -2.05740092045291e-07 wetab = -9.11009369437662e-07 petab = 6.16565152786814e-13
+ dsub = -0.822371491891293 ldsub = 7.58251135344101e-07 wdsub = 3.63705449519155e-06 pdsub = -2.51153508543482e-12
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 4.24164187899261 lpclm = -2.36485780726675e-06 wpclm = -6.78910421731446e-06 ppclm = 5.02900470171464e-12
+ pdiblc1 = 0.235754794952707 lpdiblc1 = 1.53483010446239e-07 wpdiblc1 = -9.94580372318717e-08 ppdiblc1 = 6.22069166350474e-14
+ pdiblc2 = -0.0481375380305695 lpdiblc2 = 4.41283817300152e-08 wpdiblc2 = 4.74827388501969e-08 ppdiblc2 = -4.26077654241674e-14
+ pdiblcb = -0.025
+ drout = 0.0655147863297549 ldrout = 1.71534022393344e-07 wdrout = 8.24252289823722e-07 pdrout = -3.2488380163007e-13
+ pscbe1 = 211361246.720848 lpscbe1 = 150.797048836316 wpscbe1 = -773.722879795036 ppscbe1 = 0.000464812868926163
+ pscbe2 = 1.61558182116595e-08 lpscbe2 = -1.80337553142229e-15 wpscbe2 = 6.03566187835619e-15 ppscbe2 = -4.17478333717877e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.000507633755157381 lalpha0 = -3.46482042890874e-10 walpha0 = -8.05289862703754e-10 palpha0 = 5.83530630966344e-16
+ alpha1 = 0.0
+ beta0 = 130.799178104221 lbeta0 = -5.99932419818279e-05 wbeta0 = -0.000193870363245486 pbeta0 = 1.37206340143981e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -8.94239537294086e-08 lagidl = 7.89134774702079e-14 wagidl = 1.77664657345649e-13 pagidl = -1.40471691685835e-19
+ bgidl = 578328462.007801 lbgidl = 854.823707501339 wbgidl = 457.573803187435 pbgidl = -0.000352654811187715
+ cgidl = 3798.2529650946 lcgidl = -0.00223864338777451 wcgidl = -0.00455568717038673 pcgidl = 3.09965018254465e-9
+ egidl = 0.185684181143102 legidl = 4.23757531527567e-07 wegidl = 4.87427766118957e-06 pegidl = -4.00771933823974e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.728600013257001 lkt1 = 6.03480685809794e-08 wkt1 = 4.06443394540008e-07 pkt1 = -2.78411693042933e-13
+ kt2 = -0.019032
+ at = 119474.287045167 lat = -0.0612426632292707 wat = -0.218530386190657 pat = 1.39205846521466e-7
+ ute = -1.70970406009967 lute = 1.57483131647971e-07 wute = 9.48367920593353e-07 pute = -6.49627283766843e-13
+ ua1 = 5.524e-10
+ ub1 = -3.5909e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.41e-6
+ sbref = 2.41e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.54 pmos
* DC IV MOS Parameters
+ lmin = 6e-07 lmax = 8.0e-07 wmin = 1.5e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.12544727723518+0*(0.0/sqrt(l*w*mult))} lvth0 = 9.50573266169239e-08 wvth0 = 3.95833343949101e-07 pvth0 = -1.46228060789218e-13
+ k1 = 0.69955473701484 lk1 = -8.48457693606602e-08 wk1 = -3.72198593007008e-07 pk1 = 2.56275458513103e-13
+ k2 = -0.0143188011413564 lk2 = 3.2973076612842e-08 wk2 = 9.58191743940365e-08 pk2 = -6.55386773646472e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 27558.0774948915 lvsat = 0.024545442583613 wvsat = -0.00178023979554687 pvsat = -6.61260867550577e-9
+ ua = 2.91264921059795e-09 lua = 2.87376385057356e-16 wua = -1.71379964335569e-15 pua = -8.68264203229374e-22
+ ub = -6.3969877188538e-19 lub = -3.44541803668348e-25 wub = 2.0273670828398e-24 pub = 5.02124945802713e-31
+ uc = -5.17346643003282e-12 luc = 1.45486466885984e-18 wuc = 8.17846854458412e-18 puc = -4.39439836418578e-24
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0264399561635315 lu0 = -2.93804950011573e-09 wu0 = -1.19305066592063e-08 pu0 = 1.43064668544823e-15
+ a0 = 1.00473103316073 la0 = -7.74539668702198e-08 wa0 = -4.8696587356753e-07 pa0 = 2.33948622575963e-13
+ keta = -0.141721898752241 lketa = 5.20261053182995e-08 wketa = 6.88137024006156e-08 pketa = -4.59353034588281e-14
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.673033935768526 lags = 2.27900215362554e-08 wags = 1.45243283806267e-07 pags = -6.88369409899588e-14
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0529144832576219+0*(0.009/sqrt(l*w*mult))} lvoff = -6.14144794921755e-09 wvoff = -6.01283549099844e-08 pvoff = 1.85501575503404e-14
+ nfactor = {1.15516476546576+0*(0.02/sqrt(l*w*mult))} lnfactor = 4.29904830648853e-07 wnfactor = 6.10432278335488e-07 pnfactor = -4.68456687510258e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.0239800182065449 leta0 = -2.01830765731097e-08 weta0 = -6.68420954788676e-08 peta0 = 5.8606367724712e-14
+ etab = 0.0105465780654758 letab = -5.11503762886541e-09 wetab = -3.73585511556898e-08 petab = 1.81187105177538e-14
+ dsub = 0.300846638333833 ldsub = -1.11476677694585e-08 wdsub = -7.85767854518823e-08 pdsub = 3.36537636495334e-14
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.659449553551769 lpclm = 8.89260246985964e-08 wpclm = 9.4466423889139e-07 ppclm = -2.68588021944089e-13
+ pdiblc1 = 0.323202059176803 lpdiblc1 = 9.35820716890546e-08 wpdiblc1 = 4.04005862537958e-07 ppdiblc1 = -2.82663337387786e-13
+ pdiblc2 = 0.0193428364891883 lpdiblc2 = -2.0953374141463e-09 wpdiblc2 = -2.39582245858464e-08 ppdiblc2 = 6.32893732470509e-15
+ pdiblcb = -0.025
+ drout = 0.552371172625675 ldrout = -1.6196016793743e-07 wdrout = -3.64197584179336e-07 pdrout = 4.89198419812656e-13
+ pscbe1 = 356779883.619084 lpscbe1 = 51.186009654208 wpscbe1 = 130.545756446926 ppscbe1 = -0.0001546066255564
+ pscbe2 = 1.63030265550921e-08 lpscbe2 = -1.90421251063191e-15 wpscbe2 = -8.45558341039378e-15 ppscbe2 = 5.75164722938853e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -5.0669632529136e-06 lalpha0 = 4.71538571658577e-12 walpha0 = 6.7378386711046e-11 palpha0 = -1.42427565415473e-17
+ alpha1 = 0.0
+ beta0 = 45.0053579977245 lbeta0 = -1.22490417797853e-06 wbeta0 = 1.03110935366493e-06 pbeta0 = 3.69980592092567e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.4672037966288e-07 lagidl = -8.28442101818427e-14 wagidl = -3.55995703144709e-13 pagidl = 2.25082986948258e-19
+ bgidl = 1236804524.81572 lbgidl = 403.770896858233 wbgidl = 1723.17359585748 pbgidl = -0.00121958434116774
+ cgidl = 1651.02729683973 lcgidl = -0.000767804541148266 wcgidl = -0.00341625211572226 pcgidl = 2.31914286727476e-9
+ egidl = 3.38797108539564 legidl = -1.7697929864509e-06 wegidl = -8.78035379847491e-06 pegidl = 5.34563493847313e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.6480883740352 lkt1 = 5.19799827224159e-09 wkt1 = 5.93971006645768e-08 pkt1 = -4.06867169697323e-14
+ kt2 = -0.019032
+ at = 39668.8305909667 lat = -0.0065763245854259 wat = 0.00696522382856346 pat = -1.52575188636497e-8
+ ute = -1.24897725987041 lute = -1.58112422875068e-07 wute = -8.6200042339469e-07 pute = 5.90465980023246e-13
+ ua1 = 5.53369990000001e-10 lua1 = -6.644383000496e-19
+ ub1 = -7.84174465559763e-19 lub1 = -1.92259295746389e-24 wub1 = -1.06142618887601e-23 pub1 = 7.27071632249123e-30
+ uc1 = -4.39803282716397e-10 luc1 = 2.26461595644319e-16 wuc1 = 5.02677662924324e-16 puc1 = -3.44331685714848e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.02e-6
+ sbref = 2.01e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.55 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 6e-07 wmin = 1.5e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.014/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.649208696256675+0*(0.0/sqrt(l*w*mult))} lvth0 = -1.35916003964743e-07 wvth0 = -1.752094654008e-07 pvth0 = 1.30724846531435e-13
+ k1 = 0.440036547081725 lk1 = 4.10192551659509e-08 wk1 = 4.99934451805871e-07 pk1 = -1.66704707555919e-13
+ k2 = 0.0773563180283725 lk2 = -1.14888978088806e-08 wk2 = -1.84939825626456e-07 pk2 = 7.06280338502914e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -198757.45676155 lvsat = 0.134307345120316 wvsat = 0.355250381698133 pvsat = -1.79770674946833e-7
+ ua = 3.84188005152506e-09 lua = -1.6329592663809e-16 wua = -7.43557104275845e-15 pua = 1.90676631662397e-21
+ ub = -6.47214514365965e-18 lub = 2.48416552441032e-24 wub = 1.39361007808825e-23 pub = -5.27355135407948e-30
+ uc = 2.54225370213859e-10 luc = -1.24352274109244e-16 wuc = -3.85372261192037e-16 puc = 1.86475737804427e-22
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.008040057040757 lu0 = 5.98580957493427e-09 wu0 = 4.1871687410357e-09 pu0 = -6.38634529529211e-15
+ a0 = 0.10373780370872 la0 = 3.5952324444786e-07 wa0 = 1.27800933586073e-06 pa0 = -6.220555291207e-13
+ keta = -0.347864105893917 lketa = 1.52004045070977e-07 wketa = 4.30914512285109e-07 pketa = -2.21552385748758e-13
+ a1 = 0.0
+ a2 = 0.5
+ ags = 5.32189917486541 lags = -2.23188637509954e-06 wags = -7.72034328016673e-06 pags = 3.74593321460413e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {0.257718857257401+0*(0.009/sqrt(l*w*mult))} lvoff = -1.56797064932301e-07 wvoff = -4.44959023439656e-07 pvoff = 2.05191107633888e-13
+ nfactor = {2.64608344218373+0*(0.02/sqrt(l*w*mult))} lnfactor = -2.93183272965978e-07 wnfactor = -2.40708863807709e-06 pnfactor = 9.95025869345259e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -0.968950598465193 leta0 = 4.613833078596e-07 weta0 = 1.258035852896e-06 peta0 = -5.83952812847356e-13
+ etab = 0.0626256364476834 letab = -3.03731205489442e-08 wetab = -1.34731552276419e-08 petab = 6.53441291963017e-15
+ dsub = 0.142824246807478 ldsub = 6.54924020088661e-08 wdsub = 1.85536885589888e-07 pdsub = -9.44400462373702e-14
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 3.43107656970022 lpclm = -1.25529921999832e-06 wpclm = -3.16481356750197e-06 ppclm = 1.72448816676766e-12
+ pdiblc1 = 1.76527724829863 lpdiblc1 = -6.05817184659088e-07 wpdiblc1 = -8.39629219221493e-07 ppdiblc1 = 3.20493459090139e-13
+ pdiblc2 = 0.0583320034843444 lpdiblc2 = -2.1004888460962e-08 wpdiblc2 = -5.35508738018298e-08 ppdiblc2 = 2.06812242312109e-14
+ pdiblcb = 1.52549601009334 lpdiblcb = -7.51982812415217e-07 wpdiblcb = -2.35750747640278e-06 ppdiblcb = 1.14337933851796e-12
+ drout = -2.79057911069841 ldrout = 1.45935400472333e-06 wdrout = 3.12564412473599e-06 pdrout = -1.20335735980273e-12
+ pscbe1 = 717713710.410581 lpscbe1 = -123.865091670534 wpscbe1 = -591.561053684649 ppscbe1 = 0.000195611566823363
+ pscbe2 = 4.84571875908612e-09 lpscbe2 = 3.65252448389199e-15 wpscbe2 = 1.40626510048406e-14 ppscbe2 = -5.16958387082804e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 9.35639499472819e-05 lalpha0 = -4.3120114030943e-11 walpha0 = -3.00549460331662e-11 palpha0 = 3.30119226727319e-17
+ alpha1 = -7.75248005046668e-10 lalpha1 = 3.75991406207609e-16 walpha1 = 1.17875373820139e-15 palpha1 = -5.71689669258982e-22
+ beta0 = 362.141459436547 lbeta0 = -0.0001550343276953 wbeta0 = -0.000464435775845631 pbeta0 = 2.29448917908158e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -2.10157615948481e-07 lagidl = 9.02398332996893e-14 wagidl = 6.16537815381089e-13 pagidl = -2.46590906869162e-19
+ bgidl = 7161306612.28024 lbgidl = -2469.58299305163 wbgidl = -9343.31758784885 pbgidl = 0.00414760855047392
+ cgidl = -3676.54126832107 lcgidl = 0.0018160395751119 wcgidl = 0.00978678750818063 pcgidl = -4.08426533512002e-9
+ egidl = -14.2653921133374 legidl = 6.79199989811865e-06 wegidl = 2.68777867150064e-05 pegidl = -1.19483849198628e-11
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.993459023150135 lkt1 = 1.7270103623974e-07 wkt1 = 3.99857443479458e-07 pkt1 = -2.05808280933235e-13
+ kt2 = -0.019032
+ at = 6596.60841433328 lat = 0.00946353780913042 wat = 0.034443784637024 pat = -2.85844834629491e-8
+ ute = -2.84607392763188 lute = 6.16471475505904e-07 wute = 2.04462186358016e-06 pute = -8.19231296048123e-13
+ ua1 = 5.52e-10
+ ub1 = -9.02292416683795e-18 lub1 = 2.07315945390752e-24 wub1 = 1.25764713391221e-23 pub1 = -3.97667333936548e-30
+ uc1 = 2.7132656096e-11 wuc1 = -2.07291894936783e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 1.81e-6
+ sbref = 1.81e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.56 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 1e-06 wmax = 1.5e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.937322024208+0*(0.0/sqrt(l*w*mult))} wvth0 = 1.10600519719248e-8
+ k1 = 0.57432823688 wk1 = 1.07373119592763e-8
+ k2 = 0.02454322024768 wk2 = -4.20306801087972e-10
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 384843.148568 wvsat = -0.310928969493564
+ ua = 3.55426774524664e-09 wua = -1.3307676106052e-15
+ ub = -8.58442672480001e-19 wub = 1.08254448088843e-24
+ uc = 2.0155487937704e-11 wuc = -6.66010696744479e-17
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.02195954085716 wu0 = -3.25542264873979e-9
+ a0 = 1.06718596410856 wa0 = -1.63927038205368e-7
+ keta = -0.0125572505136 wketa = 4.46498394422161e-9
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.17929876938976 wags = -5.42950488509986e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.081326978459812+0*(0.009/sqrt(l*w*mult))} wvoff = -2.68930222026404e-8
+ nfactor = {1.65144+0*(0.02/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 5.0e-6
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.0800000000000101
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.38907759208228 wpclm = -2.35277776444618e-6
+ pdiblc1 = 0.39
+ pdiblc2 = -0.0030941437847352 wpdiblc2 = 6.66602924667689e-9
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 205246692.02008 wpscbe1 = 19.8697992056567
+ pscbe2 = 1.495748741968e-08 wpscbe2 = 4.20803324184346e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -6.98392547789081e-05 walpha0 = 1.36828697495835e-10
+ alpha1 = 0.0
+ beta0 = 34.264470782272 wbeta0 = 4.8728280155904e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -1.10179144e-08 wagidl = 3.16533473943984e-14
+ bgidl = 2348456675.6 wbgidl = -845.020244656343
+ cgidl = -1434.185904 wcgidl = 0.00289224703642935
+ egidl = -0.389880758542361 wegidl = 1.94894044826906e-6
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.67763888 wkt1 = 1.24130774095679e-7
+ kt2 = -0.019032
+ at = 730334.34656 wat = -0.591110746243629
+ ute = -1.5561
+ ua1 = 2.2096e-11
+ ub1 = -5.1351339468e-18 wub1 = 2.10060302463415e-24
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.57 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 1e-06 wmax = 1.5e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.937322024208+0*(0.0/sqrt(l*w*mult))} wvth0 = 1.10600519719252e-8
+ k1 = 0.57432823688 wk1 = 1.07373119592768e-8
+ k2 = 0.02454322024768 wk2 = -4.20306801087972e-10
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 384843.148568 wvsat = -0.310928969493564
+ ua = 3.55426774524664e-09 wua = -1.3307676106052e-15
+ ub = -8.58442672480001e-19 wub = 1.08254448088843e-24
+ uc = 2.0155487937704e-11 wuc = -6.66010696744479e-17
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.02195954085716 wu0 = -3.25542264873978e-9
+ a0 = 1.06718596410856 wa0 = -1.63927038205368e-7
+ keta = -0.0125572505136 wketa = 4.46498394422161e-9
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.17929876938976 wags = -5.42950488509986e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.081326978459812+0*(0.009/sqrt(l*w*mult))} wvoff = -2.68930222026404e-8
+ nfactor = {1.65144+0*(0.02/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 5.0e-6
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.0800000000000101
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.38907759208228 wpclm = -2.35277776444618e-6
+ pdiblc1 = 0.39
+ pdiblc2 = -0.0030941437847352 wpdiblc2 = 6.66602924667689e-9
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 205246692.02008 wpscbe1 = 19.8697992056566
+ pscbe2 = 1.495748741968e-08 wpscbe2 = 4.20803324184219e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -6.98392547789081e-05 walpha0 = 1.36828697495835e-10
+ alpha1 = 0.0
+ beta0 = 34.264470782272 wbeta0 = 4.8728280155904e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -1.10179144e-08 wagidl = 3.16533473943984e-14
+ bgidl = 2348456675.6 wbgidl = -845.020244656343
+ cgidl = -1434.185904 wcgidl = 0.00289224703642935
+ egidl = -0.389880758542361 wegidl = 1.94894044826906e-6
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.677638879999999 wkt1 = 1.2413077409568e-7
+ kt2 = -0.019032
+ at = 730334.34656 wat = -0.591110746243629
+ ute = -1.5561
+ ua1 = 2.2096e-11
+ ub1 = -5.1351339468e-18 wub1 = 2.10060302463415e-24
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.58 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 1e-06 wmax = 1.5e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.905559767442853+0*(0.0/sqrt(l*w*mult))} lvth0 = -2.504452357819e-07 wvth0 = -3.72340147678872e-08 pvth0 = 3.8079847477308e-13
+ k1 = 0.614469639831646 lk1 = -3.16514761566716e-07 wk1 = -5.0297129249061e-08 pk1 = 4.81256263755532e-13
+ k2 = 0.0124290721264132 lk2 = 9.55199973654485e-08 wk2 = 1.79990858192246e-08 pk2 = -1.45236818714201e-13
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 464281.49829068 lvsat = -0.626370990371585 wvsat = -0.431713868110004 pvsat = 9.5238832166613e-7
+ ua = 2.99160966465642e-09 lua = 4.43655615216347e-15 wua = -4.75253876280904e-16 pua = -6.74572151757844e-21
+ ub = -5.99535579170641e-19 lub = -2.04148113620883e-24 wub = 6.88879870210852e-25 pub = 3.10404348686962e-30
+ uc = 5.02992433358408e-11 luc = -2.37683360595531e-16 wuc = -1.12434227744739e-16 puc = 3.61394222218457e-22
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0205742560855699 lu0 = 1.09229634975639e-08 wu0 = -1.14911654752385e-09 pu0 = -1.66082130765568e-14
+ a0 = 0.992549477678819 la0 = 5.88508322316082e-07 wa0 = -5.04433054997556e-08 pa0 = -8.94818664965088e-13
+ keta = -0.0158187147247775 lketa = 2.57166289978132e-08 wketa = 9.42399461681799e-09 pketa = -3.91017743583691e-14
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.170836386783017 lags = 6.67258445422572e-08 wags = -4.14281145708021e-08 pags = -1.01455712464678e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.060295561388971+0*(0.009/sqrt(l*w*mult))} lvoff = -1.65832618446496e-07 wvoff = -5.88709974190151e-08 pvoff = 2.5214617469124e-13
+ nfactor = {1.76898988617445+0*(0.02/sqrt(l*w*mult))} lnfactor = -9.26880264736114e-07 wnfactor = -1.78732956229846e-07 pnfactor = 1.40930846620755e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.4911457518925e-05 lcit = -7.81517929794362e-11 wcit = -1.50702323971202e-11 pcit = 1.18828707100131e-16
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.0800000000000101
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 4.03456016662566 lpclm = -1.29746218728617e-05 wpclm = -4.85471098228334e-06 ppclm = 1.97277309129799e-11
+ pdiblc1 = 0.39
+ pdiblc2 = -0.00735223795547955 lpdiblc2 = 3.35750512458483e-08 wpdiblc2 = 1.31404018199753e-08 ppdiblc2 = -5.10503953685948e-14
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 205922772.360361 lpscbe1 = -5.33089010271306 wpscbe1 = 18.8418285133844 ppscbe1 = 8.10554376871366e-6
+ pscbe2 = 1.49746659578518e-08 lpscbe2 = -1.35452687591989e-16 wpscbe2 = 1.59606056277316e-17 ppscbe2 = 2.05953915146043e-22
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -0.000197186697984768 lalpha0 = 1.00413395294099e-09 walpha0 = 3.3045870202614e-10 palpha0 = -1.52677161757143e-15
+ alpha1 = 1.982291503785e-10 lalpha1 = -1.56303585958872e-15 walpha1 = -3.01404647942405e-16 palpha1 = 2.37657414200262e-21
+ beta0 = -37.1762802579746 lbeta0 = 0.000563309964748589 wbeta0 = 0.000113497489801771 pbeta0 = -8.56504915060723e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.59412500514761e-08 lagidl = -2.12572876904066e-13 wagidl = -9.33768472576862e-15 pagidl = 3.23214083312356e-19
+ bgidl = 2253108454.26794 lbgidl = 751.820248462172 wbgidl = -700.044608996046 pbgidl = -0.00114313216230326
+ cgidl = -3234.10658943679 lcgidl = 0.0141923656050656 wcgidl = 0.00562900123974638 pcgidl = -2.15792932093838e-8
+ egidl = 0.561747615763887 legidl = -7.50358497326289e-06 wegidl = 5.02002827933651e-07 pegidl = 1.14090959016566e-11
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.7172847100757 lkt1 = 3.12607171917742e-07 wkt1 = 1.8441170368416e-07 pkt1 = -4.75314828400522e-13
+ kt2 = -0.019032
+ at = 866240.2520595 lat = -1.07161738533403 wat = -0.797753772872941 pat = 1.629379231757e-6
+ ute = -1.26728012789853 lute = -2.27734324742077e-06 wute = -4.39146572052083e-07 pute = 3.46266852489781e-12
+ ua1 = 2.2096e-11
+ ub1 = -3.79332082788793e-18 lub1 = -1.05801897335561e-23 wub1 = 6.03949627120112e-26 pub1 = 1.60870303672157e-29
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.59 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 1e-06 wmax = 1.5e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.957974109261406+0*(0.0/sqrt(l*w*mult))} lvth0 = -4.6815779888534e-08 wvth0 = 3.58262169714121e-08 pvth0 = 9.69598397670629e-14
+ k1 = 0.510646193972037 lk1 = 8.6838806480638e-08 wk1 = 1.07564966652234e-07 pk1 = -1.3203718951052e-13
+ k2 = 0.0551796508277497 lk2 = -7.05657871363505e-08 wk2 = -4.40375813369747e-08 pk2 = 9.5775323004297e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 112300.274685329 lvsat = 0.74107430342909 wvsat = 0.103468654644804 pvsat = -1.12679310332368e-6
+ ua = 3.52799129450922e-09 lua = 2.35271620209349e-15 wua = -1.29021421405802e-15 pua = -3.57960468011603e-21
+ ub = -9.37818288374534e-19 lub = -7.27254502365253e-25 wub = 1.10903933749615e-24 pub = 1.47172605726356e-30
+ uc = 6.00097074730491e-11 luc = -2.75408465216265e-16 wuc = -1.08666594908919e-16 puc = 3.4675698748946e-22
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0213411061766783 lu0 = 7.94375472785823e-09 wu0 = -2.54883252394523e-09 pu0 = -1.11703235067398e-14
+ a0 = 1.5849667928591 la0 = -1.71302998507276e-06 wa0 = -8.11760475559314e-07 pa0 = 2.06289473413045e-12
+ keta = -0.21127996173805 lketa = 7.85082596338141e-07 wketa = 3.0662008424304e-07 pketa = -1.1937070965758e-12
+ a1 = 0.0
+ a2 = 0.5
+ ags = 1.3562540481727 lags = -4.53861584286836e-06 wags = -1.82672588290088e-06 pags = 6.83441719100883e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0819888793021806+0*(0.009/sqrt(l*w*mult))} lvoff = -8.15541868202661e-08 wvoff = -2.58866112384306e-08 pvoff = 1.24001999301599e-13
+ nfactor = {1.85152261654239+0*(0.02/sqrt(l*w*mult))} lnfactor = -1.24751950955192e-06 wnfactor = -1.78157034590613e-07 pnfactor = 1.40707101351873e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -1.10796072587833e-05 lcit = 2.2823363726637e-11 wcit = 2.44488177224785e-11 pcit = -3.47026050192594e-17
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -0.07388888060559 leta0 = 5.97857531708353e-07 weta0 = 2.33985888516486e-07 peta0 = -9.09034006957108e-13
+ etab = 0.0634062705969947 letab = -5.18282694237972e-07 wetab = -2.02842366754942e-07 petab = 7.88041580631117e-13
+ dsub = -0.0170833022710006 ldsub = 2.24196574390633e-06 wdsub = 8.77447081936825e-07 pdsub = -3.40887752608916e-12
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.59909130559201 lpclm = -7.39783252509023e-06 wpclm = -2.67210067564573e-06 ppclm = 1.12483007847443e-11
+ pdiblc1 = 0.391747215878176 lpdiblc1 = -6.78792495063387e-09 wpdiblc1 = -2.65661728174397e-09 ppdiblc1 = 1.03209448564888e-14
+ pdiblc2 = 0.00129
+ pdiblcb = -0.025
+ drout = 0.710041985604331 ldrout = -5.82912363862899e-07 wdrout = -2.28136738523587e-07 pdrout = 8.86310088480444e-13
+ pscbe1 = 367757084.949938 lpscbe1 = -634.056385341657 wpscbe1 = -227.224978098691 ppscbe1 = 0.000964073857122594
+ pscbe2 = 1.44791378394572e-08 lpscbe2 = 1.78967157473066e-15 wpscbe2 = 7.69404172253168e-16 ppscbe2 = -2.72117057397595e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.000676385851515773 lalpha0 = -2.38969103400587e-09 walpha0 = -9.9779612947374e-10 palpha0 = 3.63349176153144e-15
+ alpha1 = -3.96458300757e-10 lalpha1 = 7.47321914635442e-16 walpha1 = 6.02809295884808e-16 palpha1 = -1.13629250869638e-21
+ beta0 = 208.508645994069 lbeta0 = -0.000391174745315968 wbeta0 = -0.000260063000975494 pbeta0 = 5.94775723806495e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -5.5698329928766e-08 lagidl = 6.57465331212743e-14 wagidl = 8.49721402914628e-14 pagidl = -4.31791153304627e-20
+ bgidl = 3253050998.71177 lbgidl = -3132.95153698936 wbgidl = -1945.44013732591 pbgidl = 0.00369522323828065
+ cgidl = -1009.55812490688 lcgidl = 0.00555000594310925 wcgidl = 0.00119761072933654 pcgidl = -4.36336323339412e-9
+ egidl = -2.41406492842354 legidl = 4.05743188184254e-06 wegidl = 5.02668413999501e-06 pegidl = -6.16926837229525e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.72903692034065 lkt1 = 3.58264450036023e-07 wkt1 = 1.93682449338364e-07 pkt1 = -5.11331628913373e-13
+ kt2 = -0.019032
+ at = 343776.116324728 lat = 0.958153169674884 wat = 0.0683986575008948 pat = -1.73561862948321e-6
+ ute = -2.26008546240753 lute = 1.57970051312004e-06 wute = 8.60744202465427e-07 pute = -1.58740063464885e-12
+ ua1 = -5.26731060073324e-11 lua1 = 2.90477602992957e-16 wua1 = -6.46269024082536e-16 pua1 = 2.51075192721553e-21
+ ub1 = -5.85718029090663e-18 lub1 = -2.56210603902575e-24 wub1 = 3.9139883711143e-24 pub1 = 1.11583924353985e-30
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.60 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 1e-06 wmax = 1.5e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.980816602436167+0*(0.0/sqrt(l*w*mult))} lvth0 = -3.7577944665761e-09 wvth0 = 6.57076143620396e-08 pvth0 = 4.06335550927164e-14
+ k1 = 0.561754086062241 lk1 = -9.49931456993578e-09 wk1 = 2.98561322395685e-08 pk1 = 1.44435748131833e-14
+ k2 = 0.0159440028423889 lk2 = 3.39321313781472e-09 wk2 = 8.55891030191731e-09 pk2 = -3.36880075255617e-15
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 631045.172378248 lvsat = -0.236757234997575 wvsat = -0.644907024641612 pvsat = 2.83891310252815e-7
+ ua = 3.48198856194386e-09 lua = 2.43943112296553e-15 wua = -1.22187351477517e-15 pua = -3.70842655656069e-21
+ ub = -1.69609789272693e-19 lub = -2.17532368212973e-24 wub = 1.63369886845974e-25 pub = 3.25430824339189e-30
+ uc = -1.62365971516217e-10 luc = 1.43768577800106e-16 wuc = 1.4400471832148e-16 puc = -1.29527174593276e-22
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0221051972382718 lu0 = 6.50344689720986e-09 wu0 = -3.06032028268255e-09 pu0 = -1.02061716389588e-14
+ a0 = 0.493026960520744 la0 = 3.45271139185893e-07 wa0 = 5.43967650795408e-07 pa0 = -4.92646005407572e-13
+ keta = 0.254784921955133 lketa = -9.34473790990891e-08 wketa = -4.02025046504072e-07 pketa = 1.42085431656858e-13
+ a1 = 0.0
+ a2 = 0.5
+ ags = -0.957651591191027 lags = -1.7691528219593e-07 wags = 1.71228708006934e-06 pags = 1.63395450874777e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.113489767915232+0*(0.009/sqrt(l*w*mult))} lvoff = -2.2175169289108e-08 wvoff = 2.20100488852729e-08 pvoff = 3.37170344517187e-14
+ nfactor = {1.27338584754394+0*(0.02/sqrt(l*w*mult))} lnfactor = -1.5773459067367e-07 wnfactor = 4.9502835518487e-07 pnfactor = 1.38119919718901e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -2.48661555813334e-06 lcit = 6.62561733587021e-12 wcit = 1.13832941435239e-11 pcit = -1.00741584005479e-17
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.314700498098676 leta0 = -1.34631504202295e-07 weta0 = -3.56858821552048e-07 peta0 = 2.0470531729853e-13
+ etab = -0.211795041646092 letab = 4.70403333685436e-10 wetab = 2.155973756923e-07 petab = -7.15241683221993e-16
+ dsub = 1.25883552266291 ldsub = -1.63134861499976e-07 wdsub = -1.06256962851164e-06 pdsub = 2.48044273022652e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -2.47352855710233 lpclm = 2.16403055298929e-06 wpclm = 5.04074982309736e-06 ppclm = -3.29038384113388e-12
+ pdiblc1 = 0.269548983200817 lpdiblc1 = 2.23555132655024e-07 wpdiblc1 = 1.83144084728922e-07 ppdiblc1 = -3.39912449430106e-13
+ pdiblc2 = 0.0025953794146917 lpdiblc2 = -2.46063366979678e-09 wpdiblc2 = -1.98481112472693e-09 ppdiblc2 = 3.74135904605463e-15
+ pdiblcb = -0.025
+ drout = 1.05466543939043 ldrout = -1.23252585113243e-06 wdrout = -7.52131875277002e-07 pdrout = 1.87403830128495e-12
+ pscbe1 = 33435821.7311149 lpscbe1 = -3.86247578049188 wpscbe1 = 281.105822127844 ppscbe1 = 5.8728403495769e-6
+ pscbe2 = 1.47972585811524e-08 lpscbe2 = 1.19001556723891e-15 wpscbe2 = 2.85706038195984e-16 ppscbe2 = -1.80940200976882e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -0.00103485487396858 lalpha0 = 8.35989177328512e-10 walpha0 = 1.60412143625506e-09 palpha0 = -1.27110984027952e-15
+ alpha1 = 0.0
+ beta0 = -8.75061291512398 lbeta0 = 1.83578714315653e-05 wbeta0 = 7.02766605663092e-05 pbeta0 = -2.79128865014951e-11
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -6.86790894590207e-08 lagidl = 9.02151999320065e-14 wagidl = 1.45331169574235e-13 pagidl = -1.56955583733341e-19
+ bgidl = 1525567120.22021 lbgidl = 123.346936547825 wbgidl = 138.208058828837 pbgidl = -0.000232443193230084
+ cgidl = 2747.41192718289 lcgidl = -0.0015318638202297 wcgidl = -0.00151314972679092 pcgidl = 7.46406672603867e-10
+ egidl = -2.71278389250281 legidl = 4.62051563553715e-06 wegidl = 5.48088214281205e-06 pegidl = -7.02542933661534e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.55360700019682 lkt1 = 2.7579927714505e-08 wkt1 = -4.18788216230382e-08 pkt1 = -6.72998109574853e-14
+ kt2 = -0.019032
+ at = 1633444.48036921 lat = -1.47286524820715 wat = -1.66161505929771 pat = 1.52544857661358e-6
+ ute = -1.5562669879841 lute = 2.53006207924249e-07 wute = 1.97134177048161e-07 pute = -3.36499054787428e-13
+ ua1 = -2.97682176465336e-10 lua1 = 7.52318475760939e-16 wua1 = 1.29253804816507e-15 pua1 = -1.14388970993585e-21
+ ub1 = -1.04249330559833e-17 lub1 = 6.04808508437993e-24 wub1 = 8.49368775314846e-24 pub1 = -7.51687119309762e-30
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.81e-6
+ sbref = 2.81e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.61 pmos
* DC IV MOS Parameters
+ lmin = 8.0e-07 lmax = 1e-06 wmin = 1e-06 wmax = 1.5e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.39031166122285+0*(0.0/sqrt(l*w*mult))} lvth0 = 3.58643285084349e-07 wvth0 = 4.93922326325249e-07 pvth0 = -3.38334323921164e-13
+ k1 = 0.462177638123583 lk1 = 7.86253439735362e-08 wk1 = 2.04330512822701e-07 pk1 = -1.39965379630985e-13
+ k2 = -0.0286248720699268 lk2 = 4.28364445908395e-08 wk2 = 2.10289603504457e-08 pk2 = -1.44047326952535e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1417215.13093906 lvsat = -0.932513717474104 wvsat = -1.43424091009945 pvsat = 9.8244785221357e-7
+ ua = 2.29078788140577e-08 lua = -1.4752384620704e-14 wua = -2.39488925388458e-14 pua = 1.64048716446467e-20
+ ub = -1.39314264181856e-17 lub = 1.0003815225375e-23 wub = 1.69944488820058e-23 pub = -1.16411125119295e-29
+ uc = 6.85039917045227e-12 luc = -5.98706417574245e-18 wuc = -1.04185945117896e-17 puc = 7.1366851476033e-24
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.076635764082971 lu0 = -4.17558321075147e-08 wu0 = -6.45726989376571e-08 pu0 = 4.42319759088004e-14
+ a0 = 1.18167332080974 la0 = -2.6417744643807e-07 wa0 = -5.6186771459451e-08 pa0 = 3.84876575158681e-14
+ keta = 0.881491624107969 lketa = -6.48079676970838e-07 wketa = -1.06852362187007e-06 pketa = 7.31933338362888e-13
+ a1 = 0.0
+ a2 = 0.5
+ ags = -7.64203850980767 lags = 5.73873371884521e-06 wags = 8.39380477650373e-06 pags = -5.74971430288118e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.326685666753292+0*(0.009/sqrt(l*w*mult))} lvoff = 1.66502135203082e-07 wvoff = 2.65979088324704e-07 pvoff = -1.82194345606981e-13
+ nfactor = {-1.09445455113262+0*(0.02/sqrt(l*w*mult))} lnfactor = 1.93779232295309e-06 wnfactor = 2.88108769457868e-06 pnfactor = -1.97353066534792e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -1.2124875e-05 lcit = 1.5155428750625e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.696011601167681 leta0 = -4.72089923862849e-07 weta0 = -5.55564777404624e-07 peta0 = 3.80559094698281e-13
+ etab = -0.920812187601989 letab = 6.27947032418925e-07 wetab = 9.50436789087925e-07 petab = -6.51044448341283e-13
+ dsub = 3.84631810604095 ldsub = -2.45304401037662e-06 wdsub = -3.46162267681005e-06 pdsub = 2.3711942255015e-12
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -4.07305286999244 lpclm = 3.57960157227547e-06 wpclm = 5.85327274279081e-06 ppclm = -4.00946256244799e-12
+ pdiblc1 = 0.755125715563156 lpdiblc1 = -2.06177847601985e-07 wpdiblc1 = -8.89154250827171e-07 ppdiblc1 = 6.09066216045358e-13
+ pdiblc2 = -0.023435776076456 lpdiblc2 = 2.05768087840915e-08 wpdiblc2 = 9.92405562363464e-09 ppdiblc2 = -6.79792848191161e-15
+ pdiblcb = -0.025
+ drout = -3.36613435203599 ldrout = 2.67985986028099e-06 wdrout = 6.04202676162089e-06 pdrout = -4.1387581215765e-12
+ pscbe1 = -1134901275.13932 lpscbe1 = 1030.11001326436 wpscbe1 = 1273.25043701804 ppscbe1 = -0.000872170183105174
+ pscbe2 = 2.52439846603042e-08 lpscbe2 = -8.05528477918006e-15 wpscbe2 = -7.78276797247787e-15 ppscbe2 = 5.33115714730748e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -0.000510420941629634 lalpha0 = 3.71867769378206e-10 walpha0 = 7.42648050995147e-10 palpha0 = -5.08710201691421e-16
+ alpha1 = 0.0
+ beta0 = -109.438743736174 lbeta0 = 0.000107466363767541 wbeta0 = 0.000171408033581929 pbeta0 = -1.17413645963453e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.20611379661103e-07 lagidl = -7.73059187869573e-14 wagidl = -1.41691126579956e-13 pagidl = 9.70577132516372e-20
+ bgidl = 1241420765.53557 lbgidl = 374.815039711961 wbgidl = -550.648761034296 pbgidl = 0.000377191648064686
+ cgidl = 2751.17274133758 lcgidl = -0.00153519212195253 wcgidl = -0.00296361634928731 pcgidl = 2.03006238118006e-9
+ egidl = 10.5433315941259 legidl = -7.11108028955181e-06 wegidl = -1.0874380223187e-05 pegidl = 7.44889608098195e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.118101009623398 lkt1 = -3.5784069641302e-07 wkt1 = -5.21811793498831e-07 pkt1 = 3.57438469487733e-13
+ kt2 = -0.019032
+ at = -204874.751514001 lat = 0.154038080413333 wat = 0.274637786052016 pat = -1.88125510256701e-7
+ ute = -0.553133470533695 lute = -6.34761939351769e-07 wute = -8.10181468853447e-07 pute = 5.54970255257268e-13
+ ua1 = 5.524e-10
+ ub1 = -3.5909e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.41e-6
+ sbref = 2.41e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.62 pmos
* DC IV MOS Parameters
+ lmin = 6e-07 lmax = 8.0e-07 wmin = 1e-06 wmax = 1.5e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.865113841775001+0*(0.0/sqrt(l*w*mult))} lvth0 = -1.11459524833352e-9
+ k1 = 0.454765509750001 lk1 = 8.37026148487987e-8
+ k2 = 0.048699979954975 lk2 = -1.01306924219581e-8
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 26387.2414625001 lvsat = 0.0201964326778948
+ ua = 1.7855098332175e-09 lua = -2.83667480673322e-16
+ ub = 6.9366903475e-19 lub = -1.43020344085769e-26
+ uc = 2.05385163854999e-13 luc = -1.43526280629336e-18
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0185934474425 lu0 = -1.99713542037529e-9
+ a0 = 0.68446115 la0 = 7.64104045057505e-8
+ keta = -0.0964641966749999 lketa = 2.18151704863916e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.7685581851245 lags = -2.24829641998568e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0924599673396749+0*(0.009/sqrt(l*w*mult))} lvoff = 6.05870223325063e-9
+ nfactor = {1.55663658325+0*(0.02/sqrt(l*w*mult))} lnfactor = 1.21808151356666e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -0.0199809886549899 leta0 = 1.83614202027317e-08 peta0 = -6.31088724176809e-30
+ etab = -0.0140235601375 letab = 6.80135654888681e-9
+ dsub = 0.249167908341 ldsub = 1.09858892968566e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.280740534785 lpclm = -8.77201410300512e-8
+ pdiblc1 = 0.5889104330375 lpdiblc1 = -9.23212101483223e-8
+ pdiblc2 = 0.00358588470808251 lpdiblc2 = 2.06710625498653e-9
+ pdiblcb = -0.025
+ drout = 0.312844084458249 ldrout = 1.59778026174621e-7
+ pscbe1 = 442637797.76425 lpscbe1 = -50.4963639792227
+ pscbe2 = 1.074192082285e-08 lpscbe2 = 1.87855643915687e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.9246754013175e-05 lalpha0 = -4.65185379863981e-12
+ alpha1 = 0.0
+ beta0 = 45.6835025868 lbeta0 = 1.20840064753492e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -8.741245888e-08 lagidl = 6.51893704945056e-14 wagidl = -1.26217744835362e-29
+ bgidl = 2370109005.0 lbgidl = -398.330760879975
+ cgidl = -595.788600000001 lcgidl = 0.000757459662057001
+ egidl = -2.38673108119775 legidl = 1.7459479927315e-06 wegidl = -4.2351647362715e-22 pegidl = 2.01948391736579e-28
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.609023824499999 lkt1 = -2.15610228366218e-8
+ kt2 = -0.019032
+ at = 44249.75 lat = -0.01661095750125
+ ute = -1.815901535 lute = 2.30227870967326e-7
+ ua1 = 5.53369989999999e-10 lua1 = -6.64438300050389e-19
+ ub1 = -7.7650094675e-18 lub1 = 2.85924411469016e-24
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.02e-6
+ sbref = 2.01e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.63 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 6e-07 wmin = 1e-06 wmax = 1.5e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.023/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.729341944507711+0*(0.0/sqrt(l*w*mult))} lvth0 = -6.69632865634831e-08 wvth0 = -5.3367983300577e-08 pvth0 = 2.58832050608628e-14
+ k1 = 0.524227324586917 lk1 = 5.00139819619679e-08 wk1 = 3.7192355328011e-07 pk1 = -1.80381063723087e-13
+ k2 = 0.00470433592727154 lk2 = 1.1206974953258e-08 wk2 = -7.44735039694811e-08 pk2 = 3.61192770576785e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 245148.574030328 lvsat = -0.0859017198108389 wvsat = -0.319702523436486 pvsat = 1.55054125354079e-7
+ ua = -5.1221972234064e-09 lua = 3.06653590325399e-15 wua = 6.194182956693e-15 pua = -3.00414776308132e-21
+ ub = 8.42422433762056e-18 lub = -3.76358270352429e-24 wub = -8.71362046623139e-24 pub = 4.22606235801989e-30
+ uc = -1.71405433566041e-11 luc = 6.9774257964867e-18 wuc = 2.72358112690613e-17 puc = -1.32092322864384e-23
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.00843471493594367 lu0 = 2.929799051642e-09 wu0 = 3.58709693661486e-09 pu0 = -1.73972407877353e-15
+ a0 = 0.200067573260908 la0 = 3.11338867256327e-07 wa0 = 1.13154126987341e-06 pa0 = -5.48791858182255e-13
+ keta = 0.246904588319301 lketa = -1.44716973391919e-07 wketa = -4.7342296050437e-07 pketa = 2.29607768729817e-13
+ a1 = 0.0
+ a2 = 0.5
+ ags = -5.49594231187121 lags = 3.01576845434058e-06 wags = 8.72803325063548e-06 pags = -4.23305248639196e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.203980241558848+0*(0.009/sqrt(l*w*mult))} lvoff = 6.01454776281787e-08 wvoff = 2.57047992523068e-07 pvoff = -1.24666991133725e-13
+ nfactor = {0.234233366231837+0*(0.02/sqrt(l*w*mult))} lnfactor = 7.63167099594388e-07 wnfactor = 1.26009563650669e-06 pnfactor = -6.11140083227563e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -2.9288200757e-05 lcit = 1.90545809261412e-11 wcit = 5.97371592162079e-11 pcit = -2.89722235340648e-17
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.621723327316855 leta0 = -2.92861964522033e-07 weta0 = -1.16056158182064e-06 peta0 = 5.62866564375104e-13
+ etab = 0.0774867673670766 letab = -3.75806947391953e-08 wetab = -3.60692967347464e-08 petab = 1.74934285698683e-14
+ dsub = 0.300756108303254 ldsub = -1.40341297438366e-08 wdsub = -5.45962987683794e-08 pdsub = 2.64789319211703e-14
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -1.74806671477358 lpclm = 1.38123623096961e-06 wpclm = 4.71000128853447e-06 ppclm = -2.28432707493277e-12
+ pdiblc1 = 0.787365938875162 lpdiblc1 = -1.8857113820206e-07 wpdiblc1 = 6.47271235998562e-07 ppdiblc1 = -3.13923313103123e-13
+ pdiblc2 = 0.00892818454670884 lpdiblc2 = -5.23882455248062e-10 wpdiblc2 = 2.15669412393799e-08 ppdiblc2 = -1.04598586663931e-14
+ pdiblcb = -1.59652803028 lpdiblcb = 7.62183237045649e-07 wpdiblcb = 2.38948636864832e-06 ppdiblcb = -1.15888894136259e-12
+ drout = -0.734891570835499 ldrout = 6.67924580313814e-7
+ pscbe1 = 3934654077.34126 lpscbe1 = -1744.10679949268 wpscbe1 = -5482.87384443762 ppscbe1 = 0.00265916640018302
+ pscbe2 = -5.71260296698522e-08 lpscbe2 = 3.4794173088365e-14 wpscbe2 = 1.08289826886563e-13 ppscbe2 = -5.25200245908487e-20
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -3.76973800755467e-05 lalpha0 = 3.26656665137198e-11 walpha0 = 1.69526068607925e-10 palpha0 = -8.22192956445004e-17
+ alpha1 = 0.0
+ beta0 = -5.18596759208413 lbeta0 = 2.58798393369429e-05 wbeta0 = 9.40804343674249e-05 pbeta0 = -4.56285402660293e-11
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 2.26192171837654e-07 lagidl = -8.69073073804029e-14 wagidl = -4.69259280507e-14 pagidl = 2.27588404749492e-20
+ bgidl = 3838816257.38288 lbgidl = -1110.64643474941 wbgidl = -4291.51751809238 pbgidl = 0.00208136453868721
+ cgidl = 1188.54866972 lcgidl = -0.000107934992070851 wcgidl = 0.00238948636864832 pcgidl = -1.15888894136259e-9
+ egidl = -0.571595769047427 legidl = 8.65616442015158e-07 wegidl = 6.05656108666229e-06 pegidl = -2.93740184422578e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.494749795457999 lkt1 = -7.69833555518476e-08 wkt1 = -3.58422955297249e-07 pkt1 = 1.73833341204389e-13
+ kt2 = -0.019032
+ at = -2180.81060560001 lat = 0.00590763223966298 wat = 0.0477897273729664 pat = -2.31777788272518e-8
+ ute = -0.882175876069681 lute = -2.22624404985586e-07 wute = -9.41457629247438e-07 pute = 4.56602242896862e-13
+ ua1 = 5.52e-10
+ ub1 = -7.51574519999999e-19 lub1 = -5.422367676726e-25
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 1.81e-6
+ sbref = 1.81e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.64 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 7.5e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.974201738951999+0*(0.0/sqrt(l*w*mult))} wvth0 = 4.86952845521709e-8
+ k1 = 0.62747328552 wk1 = -4.34964661471628e-8
+ k2 = 0.011398456543144 wk2 = 1.29937405326992e-8
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -228636.297136 wvsat = 0.315118216135128
+ ua = 1.99244264317312e-09 wua = 2.63053040509396e-16
+ ub = 5.96488998719999e-19 wub = -4.02192920527778e-25
+ uc = -8.35391354274079e-11 wuc = 3.92178417449218e-17
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.016023457896 wu0 = 2.80226690796254e-9
+ a0 = 0.99860652433568 wa0 = -9.39426800293004e-8
+ keta = -0.0096741772848 wketa = 1.52284807725641e-9
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.13131350691392 wags = -5.32676028807861e-9
+ b0 = -1.959345898e-07 wb0 = 1.99948505806643e-13
+ b1 = -6.36575533199999e-10 wb1 = 6.49616419573135e-16
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.10350837978216+0*(0.009/sqrt(l*w*mult))} wvoff = -4.25721269280266e-9
+ nfactor = {1.3507963628+0*(0.02/sqrt(l*w*mult))} wnfactor = 3.06802622751679e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -1.040972e-05 wcit = 1.572540352392e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.0800000000000101
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -2.72541029805 wpclm = 2.86648552460335e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0100582875694704 wpdiblc2 = -6.75584281625096e-9
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 221997054.75344 wpscbe1 = 2.77628854134093
+ pscbe2 = 1.5012095555016e-08 wpscbe2 = -1.36465051780589e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.000203743717232672 walpha0 = -1.42358895280374e-10
+ alpha1 = 0.0
+ beta0 = 43.209246527848 wbeta0 = -4.25519040590951e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -1.32849951999999e-08 wagidl = 3.39668716116672e-14
+ bgidl = 961027163.999999 wbgidl = 570.832147918296
+ cgidl = 2016.3888 wcgidl = -0.0006290161409568
+ egidl = 2.8478111132304 wegidl = -1.35507877918884e-6
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.52518056 wkt1 = -3.14508070478396e-8
+ kt2 = -0.019032
+ at = -466377.480399999 wat = 0.630116919203474
+ ute = -2.0051392408 wute = 4.58238258687028e-7
+ ua1 = 2.2096e-11
+ ub1 = -5.1628678936e-18 wub1 = 2.12890512906829e-24
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.65 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 7.5e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.00555625003932+0*(0.0/sqrt(l*w*mult))} lvth0 = 6.23484296198776e-07 wvth0 = 8.06921241536244e-08 pvth0 = -6.3625699549071e-13
+ k1 = 0.655480318287397 lk1 = -5.56919706544544e-07 wk1 = -7.20772509878331e-08 pk1 = 5.68328763652811e-13
+ k2 = 0.00303188911582425 lk2 = 1.66369151459417e-07 wk2 = 2.1531705460335e-08 pk2 = -1.69777389896214e-13
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -431538.440382322 lvsat = 4.03470810394241 wvsat = 0.522177012687995 pvsat = -4.11736313415978e-6
+ ua = 1.82306485739659e-09 lua = 3.36807642327737e-15 wua = 4.35900699605343e-16 pua = -3.43707483688463e-21
+ ub = 8.55457859912683e-19 lub = -5.14959450997221e-24 wub = -6.66467017810855e-25 pub = 5.2550891031035e-30
+ uc = -1.08791195562603e-10 luc = 5.0213708952806e-16 wuc = 6.49872155840469e-17 puc = -5.12423869944132e-22
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0142191002535017 lu0 = 3.58796426992901e-08 wu0 = 4.64358862112504e-09 pu0 = -3.66146730596279e-14
+ a0 = 1.05909547782758 la0 = -1.20282253774169e-06 wa0 = -1.55670810222437e-07 pa0 = 1.22746356024987e-12
+ keta = -0.0106547271955718 lketa = 1.94982300729477e-08 wketa = 2.52348553350029e-09 pketa = -1.98976708142221e-14
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.134743366007014 lags = -6.82027309168733e-08 wags = -8.82688347455352e-09 pags = 6.9599932062437e-14
+ b0 = -3.24679861541671e-07 lb0 = 2.56009908485677e-12 wb0 = 3.31331253185213e-13 pb0 = -2.61254527470914e-18
+ b1 = -1.05485844123369e-09 lb1 = 8.31755353483547e-15 wb1 = 1.07646827126081e-15 pb1 = -8.48794693655011e-21
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.100767193981417+0*(0.009/sqrt(l*w*mult))} lvoff = -5.45084659418479e-08 wvoff = -7.0545544258599e-09 pvoff = 5.56251263751327e-14
+ nfactor = {1.15324856479135+0*(0.02/sqrt(l*w*mult))} lnfactor = 3.92823697566303e-06 wnfactor = 5.08397384950335e-07 pnfactor = -4.00871083834646e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -2.05351837626166e-05 lcit = 2.01344796292313e-10 wcit = 2.60582975371776e-11 pcit = -2.05469545789158e-16
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.0800000000000101
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -4.57111780318887 lpclm = 3.6701884511149e-05 wpclm = 4.7500041936925e-06 ppclm = -3.74537593172444e-11
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0144083216730678 lpdiblc2 = -8.65004063998645e-08 wpdiblc2 = -1.11949917184947e-08 ppdiblc2 = 8.82724537253721e-14
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 220209424.377078 lpscbe1 = 35.5470210958156 wpscbe1 = 4.60054031359368 ppscbe1 = -3.62752373699836e-5
+ pscbe2 = 1.50208824324692e-08 lpscbe2 = -1.74727014222545e-16 wpscbe2 = -2.26133906027599e-17 ppscbe2 = 1.78306471835809e-22
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.000295407491281775 lalpha0 = -1.82273368864754e-09 walpha0 = -2.35900493404647e-10 palpha0 = 1.86007421099318e-15
+ alpha1 = 0.0
+ beta0 = 45.9491301939512 lbeta0 = -5.44825730010444e-05 wbeta0 = -7.05120332879653e-06 pbeta0 = 5.55987029915439e-11
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -3.51559969272519e-08 lagidl = 4.34904759991397e-13 wagidl = 5.62859226803036e-14 pagidl = -4.43814218904581e-19
+ bgidl = 593472829.417017 lbgidl = 7308.81610541098 wbgidl = 945.916200599548 pbgidl = -0.00745854451214643
+ cgidl = 2421.40735050467 lcgidl = -0.00805379185169253 wcgidl = -0.0010423319014871 pcgidl = 8.21878183156631e-9
+ egidl = 3.72033569126724 legidl = -1.73501468716398e-05 wegidl = -2.24547789573134e-06 pegidl = 1.77055819804522e-11
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.504929632474767 lkt1 = -4.02689592584621e-07 wkt1 = -5.21165950743547e-08 pkt1 = 4.1093909157831e-13
+ kt2 = -0.019032
+ at = -872104.813368049 lat = 8.067885987433 wat = 1.04415598231471 pat = -8.23316469977156e-6
+ ute = -2.30019525484265 lute = 5.86718736395801e-06 wute = 7.59338790233354e-07 pute = -5.98738256429606e-12
+ ua1 = 2.2096e-11
+ ub1 = -6.53365317778304e-18 lub1 = 2.72580585220534e-23 wub1 = 3.5277723205831e-24 pub1 = -2.78164671089362e-29
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.66 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 7.5e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.943662719220338+0*(0.0/sqrt(l*w*mult))} lvth0 = 1.35454115158767e-07 wvth0 = 1.64951407971253e-09 pvth0 = -1.30064102709584e-14
+ k1 = 0.463169381314515 lk1 = 9.59451069931961e-07 wk1 = 1.04102666364053e-07 pk1 = -8.20849003767228e-13
+ k2 = 0.0607264550676369 lk2 = -2.88552212597797e-07 wk2 = -3.12877173089332e-08 pk2 = 2.46703494542352e-13
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 221193.433157608 lvsat = -1.11207945526058 wvsat = -0.183645900874615 pvsat = 1.44804701016684e-6
+ ua = 3.62589216168315e-09 lua = -1.08472078568856e-14 wua = -1.12253028454172e-15 pua = 8.85114568096002e-21
+ ub = -6.98231771476769e-19 lub = 7.10124046508547e-24 wub = 7.89597952712562e-25 pub = -6.2259759091488e-30
+ uc = -6.80704658180951e-11 luc = 1.81054339096261e-16 wuc = 8.36040327092426e-18 puc = -6.59217379892215e-23
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.024207100366675 lu0 = -4.28756882530807e-08 wu0 = -4.85638327657168e-09 pu0 = 3.82925578538513e-14
+ a0 = 0.966412636719459 la0 = -4.7201879901835e-07 wa0 = -2.37710252165024e-08 pa0 = 1.87434414977004e-13
+ keta = -0.00020959913012969 lketa = -6.2861552497423e-08 wketa = -6.50488931990174e-09 pketa = 5.12910197629787e-14
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.137948694848125 lags = -9.34767328023925e-08 wags = -7.86668537893218e-09 pags = 6.20287748794538e-14
+ b0 = 1.90301225425013e-07 lb0 = -1.5005242109701e-12 wb0 = -1.94199736329069e-13 pb0 = 1.53126394995603e-18
+ b1 = 6.18273190901083e-10 lb1 = -4.87508101888909e-15 wb1 = -6.30939135489882e-16 pb1 = 4.97495192864205e-21
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.153794771326071+0*(0.009/sqrt(l*w*mult))} lvoff = 3.63613716282866e-07 wvoff = 3.65436373328567e-08 pvoff = -2.88146397651389e-13
+ nfactor = {1.70833998447705+0*(0.02/sqrt(l*w*mult))} lnfactor = -4.48656093101641e-07 wnfactor = -1.16840580646276e-07 pnfactor = 9.21287394192974e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.43756250000002e-07 lcit = 3.82914576875313e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.0800000000000101
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.479252931720122 lpclm = 4.43755045894226e-06 wpclm = -2.48427908804847e-07 ppclm = 1.95885281878667e-12
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00552437360016675 lpdiblc2 = -1.64505202647798e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 226007785.201966 lpscbe1 = -10.1730250166211 wpscbe1 = -1.65464590129341 ppscbe1 = 1.30468746584698e-5
+ pscbe2 = 1.49513778463128e-08 lpscbe2 = 3.73316300097846e-16 wpscbe2 = 3.97257974197412e-17 ppscbe2 = -3.13237714025696e-22
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.000183447281497082 lalpha0 = -9.39927994296286e-10 walpha0 = -5.79729451593751e-11 palpha0 = 4.57116382716947e-16
+ alpha1 = -3.96458300757e-10 lalpha1 = 3.12607171917744e-15 walpha1 = 3.05465570317058e-16 palpha1 = -2.40859449462215e-21
+ beta0 = 177.871097610031 lbeta0 = -0.001094686626467 wbeta0 = -0.000105955348649239 pbeta0 = 8.35457394322506e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -1.59031892119602e-09 lagidl = 1.70239556742036e-13 wagidl = 8.55303596887761e-15 pagidl = -6.74406458494203e-20
+ bgidl = 2254386610.41307 lbgidl = -5787.48075317402 wbgidl = -701.348949447964 pbgidl = 0.00553013295965245
+ cgidl = 4401.17451935956 lcgidl = -0.0236642460792775 wcgidl = -0.00216269623784477 pcgidl = 1.70528490219248e-8
+ egidl = -1.67301936949262 legidl = 2.51764308156765e-05 wegidl = 2.78255124965013e-06 pegidl = -2.1940402690735e-11
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.5066416824243 lkt1 = -3.89190087292809e-07 wkt1 = -3.05465570317059e-08 pkt1 = 2.40859449462215e-13
+ kt2 = -0.019032
+ at = 478992.70750515 lat = -2.58551120916457 wat = -0.40257307512085 pat = 3.17428668446253e-6
+ ute = -1.697610942875 lute = 1.11581307701466e-6
+ ua1 = 2.2096e-11
+ ub1 = -3.734138278875e-18 lub1 = 5.18389754173799e-24
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.67 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 7.5e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.87358569585581+0*(0.0/sqrt(l*w*mult))} lvth0 = -1.36794770227305e-07 wvth0 = -5.02909774712103e-08 pvth0 = 1.88782139701914e-13
+ k1 = 0.722362551256662 lk1 = -4.75130993274318e-08 wk1 = -1.08488611927724e-07 pk1 = 5.06704943993411e-15
+ k2 = -0.0187801054828894 lk2 = 2.03303776081954e-08 wk2 = 3.14373145414443e-08 pk2 = 3.01705942879437e-15
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -96457.1391978074 lvsat = 0.121991430087354 wvsat = 0.31650267290875 pvsat = -4.95027698238668e-7
+ ua = 1.16727418264113e-09 lua = -1.29548930139725e-15 wua = 1.11886454856381e-15 pua = 1.43337961319221e-22
+ ub = -5.7759942080926e-19 lub = 6.63258438590396e-24 wub = 7.4144102620994e-25 pub = -6.03888649047074e-30
+ uc = -2.43576524403575e-12 luc = -7.39361444604571e-17 wuc = -4.49418642377519e-17 puc = 1.41157304770648e-22
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0101300028851874 lu0 = 1.18137650770114e-08 wu0 = 8.89194142957518e-09 pu0 = -1.51196148879056e-14
+ a0 = 0.121890257243882 la0 = 2.80894642263237e-06 wa0 = 6.81288645964522e-07 pa0 = -2.55171888226293e-12
+ keta = 0.30210714307075 lketa = -1.23736058436413e-06 wketa = -2.17284268794873e-07 pketa = 8.70167855126346e-13
+ a1 = 0.0
+ a2 = 0.5
+ ags = -1.25942561380097 lags = 5.33531546942782e-06 wags = 8.42538592627991e-07 pags = -3.24179147815106e-12
+ b0 = -1.05713846359752e-07 lb0 = -3.50507137161647e-13 wb0 = 1.07879500216277e-13 pb0 = 3.57687626373541e-19
+ b1 = -1.05059172779193e-09 lb1 = 1.60845084590869e-15 wb1 = 1.07211414992748e-15 pb1 = -1.64140156993798e-21
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.00545834972912762+0*(0.009/sqrt(l*w*mult))} lvoff = -2.12672539939153e-07 wvoff = -1.03984945240317e-07 pvoff = 2.57806443002479e-13
+ nfactor = {1.97027953125837+0*(0.02/sqrt(l*w*mult))} lnfactor = -1.46628992264932e-06 wnfactor = -2.99346803461459e-07 pnfactor = 1.63032315729884e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 2.17494945175667e-05 lcit = -4.56467274532739e-11 wcit = -9.05282103286186e-12 pcit = 3.51701644485632e-17
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.329683270908409 leta0 = -9.70018259062779e-07 weta0 = -1.77853842093429e-07 peta0 = 6.90961287263762e-13
+ etab = -0.133481825134189 letab = 2.466265732372e-07 wetab = -1.92082149460903e-09 petab = 7.46238190244862e-15
+ dsub = 1.00528517259906 ldsub = -1.7299306691215e-06 wdsub = -1.65865633509429e-07 pdsub = 6.44387156855963e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -2.63475868900759 lpclm = 1.28116795484753e-05 wpclm = 2.66896996994324e-06 ppclm = -9.37522335316024e-12
+ pdiblc1 = 0.841442998954461 lpdiblc1 = -1.75385379372309e-06 wpdiblc1 = -4.61564868170131e-07 ppdiblc1 = 1.79317720501662e-12
+ pdiblc2 = 0.0034413975738712 lpdiblc2 = -8.35816881750177e-09 wpdiblc2 = -2.19547110456953e-09 ppdiblc2 = 8.52939426389712e-15
+ pdiblcb = -0.025
+ drout = -0.129777367931334 ldrout = 2.6797816255264e-06 wdrout = 6.28887154288611e-07 pdrout = -2.44322344997548e-12
+ pscbe1 = 49579456.9660234 lpscbe1 = 675.250148038374 wpscbe1 = 97.4708367721023 ppscbe1 = -0.00037205512990026
+ pscbe2 = 1.45733156780717e-08 lpscbe2 = 1.84208593340364e-15 wpscbe2 = 6.73297006436744e-16 ppscbe2 = -2.77465869320066e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -0.00134383396351767 lalpha0 = 4.9935520061798e-09 walpha0 = 1.06380990869048e-09 palpha0 = -3.90100439557547e-15
+ alpha1 = 1.083389053028e-09 lalpha1 = -2.62312785104051e-15 walpha1 = -9.0735421078983e-16 palpha1 = 2.30320429087921e-21
+ beta0 = -406.033862742117 lbeta0 = 0.0011737812249763 wbeta0 = 0.000367069025594663 pbeta0 = -1.00223993449318e-9
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -7.15515538544089e-08 lagidl = 4.42038604651394e-13 wagidl = 1.01150133362446e-13 pagidl = -4.27179906237948e-19
+ bgidl = -1704190525.51343 lbgidl = 9591.57162701478 wbgidl = 3113.35543676456 pbgidl = -0.00928997450726128
+ cgidl = -1663.62909115292 lcgidl = -0.000102514376454598 wcgidl = 0.0018650809933971 pcgidl = 1.40495461743632e-9
+ egidl = 6.37505868752733 legidl = -6.09031219545577e-06 wegidl = -3.94249346235223e-06 pegidl = 4.1863623901706e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.69496519165102 lkt1 = 3.42445804435454e-07 wkt1 = 1.58912727214798e-07 pkt1 = -4.9518892253903e-13
+ kt2 = -0.019032
+ at = -326000.884455324 lat = 0.541884870633914 wat = 0.751896709918928 pat = -1.31082265806808e-6
+ ute = -1.55023781119644 lute = 5.43269197309112e-07 wute = 1.3635461227163e-07 pute = -5.29736986902216e-13
+ ua1 = -1.32779637070533e-09 lua1 = 5.24432511072837e-15 wua1 = 6.54976415816069e-16 pua1 = -2.54458010056335e-21
+ ub1 = -4.3164966197106e-18 lub1 = 7.44635678409257e-24 wub1 = 2.34174225423015e-24 pub1 = -9.09765694897287e-30
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.68 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 7.5e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.962144024357118+0*(0.0/sqrt(l*w*mult))} lvth0 = 3.01372362060161e-08 wvth0 = 4.66525098484639e-08 pvth0 = 6.04415082176538e-15
+ k1 = 0.687077721075519 lk1 = 1.89986291398707e-08 wk1 = -9.80348827605922e-08 pk1 = -1.46381777714628e-14
+ k2 = -0.00966825959626094 lk2 = 3.15459367113008e-09 wk2 = 3.46958655488853e-08 pk2 = -3.12529292747702e-15
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -36020.0266594827 lvsat = 0.00806777513817425 wvsat = 0.0358236720636053 pvsat = 3.4050814959425e-8
+ ua = 3.06601450466137e-09 lua = -4.8746053147038e-15 wua = -7.97377812955192e-16 pua = 3.75544523157073e-21
+ ub = 8.33702762145071e-19 lub = 3.97228682754596e-24 wub = -8.60496525500134e-25 pub = -3.01924221518501e-30
+ uc = -7.81297217940694e-11 luc = 6.87465851665736e-17 wuc = 5.80428047875243e-17 puc = -5.29682814186527e-23
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0232473891144075 lu0 = -1.29124423781374e-08 wu0 = -4.2259111015928e-09 pu0 = 9.6074715440833e-15
+ a0 = 1.90977456955752 la0 = -5.61206566657269e-07 wa0 = -9.01803449760093e-07 pa0 = 4.32401802717493e-13
+ keta = -0.441011471661776 lketa = 1.63414288813606e-07 wketa = 3.08025432032473e-07 pketa = -1.20038304384697e-13
+ a1 = 0.0
+ a2 = 0.5
+ ags = 1.60736816580942 lags = -6.85764711688733e-08 wags = -9.05279671673015e-07 pags = 5.2837210965021e-14
+ b0 = -9.85933268716301e-08 lb0 = -3.63929280794159e-13 wb0 = 1.00613109765922e-13 pb0 = 3.71384736040508e-19
+ b1 = 2.38069916951354e-10 lb1 = -8.20669911124182e-16 wb1 = -2.42947017270019e-16 pb1 = 8.37482154923473e-22
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.141810371096489+0*(0.009/sqrt(l*w*mult))} lvoff = 4.4350338578216e-08 wvoff = 5.09108279433012e-08 pvoff = -3.41713149697753e-14
+ nfactor = {1.06763346080297+0*(0.02/sqrt(l*w*mult))} lnfactor = 2.35193406928751e-07 wnfactor = 7.04995785320609e-07 pnfactor = -2.62857600842404e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 4.56351111626666e-06 lcit = -1.32512346717404e-11 wcit = 4.18873857407217e-12 pcit = 1.02098907972906e-17
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -0.39291948386568 leta0 = 3.92084320672607e-07 weta0 = 3.6525746336283e-07 peta0 = -3.32800807964759e-13
+ etab = -0.0139852777927529 letab = 2.13761789813288e-08 wetab = 1.37352810166611e-08 petab = -2.2049293050783e-14
+ dsub = -0.0855402100260632 ldsub = 3.26269722999951e-07 wdsub = 3.09346985437201e-07 pdsub = -2.5138625379534e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 6.45797809884569 lpclm = -4.3280838329442e-06 wpclm = -4.07372767820442e-06 ppclm = 3.33472800010985e-12
+ pdiblc1 = 0.148208519068286 lpdiblc1 = -4.47110265310047e-07 wpdiblc1 = 3.06970329609674e-07 ppdiblc1 = 3.44492199877677e-13
+ pdiblc2 = -0.00360341482992579 lpdiblc2 = 4.92126733959356e-09 wpdiblc2 = 4.34097161878581e-09 ppdiblc2 = -3.79176758741408e-15
+ pdiblcb = -0.025
+ drout = -0.0158619871151844 ldrout = 2.46505170226486e-06 wdrout = 3.4032637608801e-07 pdrout = -1.89928782587124e-12
+ pscbe1 = 403705168.958569 lpscbe1 = 7.72495156098375 wpscbe1 = -96.7488629469121 ppscbe1 = -5.95196702841603e-6
+ pscbe2 = 1.68131715227193e-08 lpscbe2 = -2.38003113447781e-15 wpscbe2 = -1.7715048958919e-15 ppscbe2 = 1.83378066867927e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.00219226579315904 lalpha0 = -1.67197835465702e-09 walpha0 = -1.68911002485934e-09 palpha0 = 1.28823591456627e-15
+ alpha1 = -3.081944e-10 walpha1 = 3.145080704784e-16
+ beta0 = 236.141298380024 lbeta0 = -3.67157428631306e-05 wbeta0 = -0.000179632106423631 pbeta0 = 2.82889658556421e-11
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 3.00655027867825e-07 lagidl = -2.59568940862109e-13 wagidl = -2.31569126480169e-13 pagidl = 1.99994234969083e-19
+ bgidl = 3610332384.29552 lbgidl = -426.277485360561 wbgidl = -1989.26570644632 pbgidl = 0.000328440834585518
+ cgidl = -1828.29350563851 lcgidl = 0.000207877221528671 wcgidl = 0.00315629360752726 pcgidl = -1.02897470413597e-9
+ egidl = 8.04653212677704 legidl = -9.24103127107428e-06 wegidl = -5.49884922443878e-06 pegidl = 7.12008521992494e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.43020834730356 lkt1 = -1.56619523375286e-07 wkt1 = -1.67805419319468e-07 pkt1 = 1.20673150087331e-13
+ kt2 = -0.019032
+ at = -99175.0165599498 lat = 0.114319243780473 wat = 0.106498880645545 pat = -9.42509768769046e-8
+ ute = -1.09585557460712 lute = -3.13239046750573e-07 wute = -2.72709224543259e-07 pute = 2.4134630017466e-13
+ ua1 = 2.25256435293067e-09 lua1 = -1.50463695152188e-15 wua1 = -1.30995283163214e-15 pua1 = 1.15930170623028e-21
+ ub1 = 2.48771078392119e-18 lub1 = -5.37954015071634e-24 wub1 = -4.68348450846031e-24 pub1 = 4.14486037256483e-30
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.81e-6
+ sbref = 2.81e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.69 pmos
* DC IV MOS Parameters
+ lmin = 8.0e-07 lmax = 1e-06 wmin = 7.5e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.04487836813388+0*(0.0/sqrt(l*w*mult))} lvth0 = 1.0335671677673e-07 wvth0 = 1.41412486794049e-07 pvth0 = -7.78179549751943e-14
+ k1 = 0.978509759203531 lk1 = -2.38917267443229e-07 wk1 = -3.22579188089692e-07 pk1 = 1.84082409723264e-13
+ k2 = -0.10372011921632 lk2 = 8.63900191755841e-08 wk2 = 9.76626087298799e-08 pk2 = -5.88505458089414e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -182157.392062778 lvsat = 0.137398612833264 wvsat = 0.197896358408614 pvsat = -1.09382702092476e-7
+ ua = -8.53849334604235e-09 lua = 5.39532611062975e-15 wua = 8.14169000132613e-15 pua = -4.15558508872917e-21
+ ub = 1.02784824920405e-17 lub = -4.38629600951284e-24 wub = -7.71142422215523e-24 pub = 3.04379454171627e-30
+ uc = -5.09122410092165e-12 luc = 4.10787990062633e-18 wuc = 1.76766485392171e-18 puc = -3.16506395311397e-24
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = -0.00316931549768601 lu0 = 1.04662091200423e-08 wu0 = 1.68672675032893e-08 pu0 = -9.05988605534433e-15
+ a0 = 2.32017275904159 la0 = -9.24406912359725e-07 wa0 = -1.21800950918292e-06 pa0 = 7.12242584276396e-13
+ keta = -0.575355864234492 lketa = 2.82308404518497e-07 wketa = 4.18168844118577e-07 pketa = -2.17514673363839e-13
+ a1 = 0.0
+ a2 = 0.5
+ ags = 1.04814587542126 lags = 4.2633245971319e-07 wags = -4.74406726041009e-07 pags = -3.28483191554578e-13
+ b0 = -2.25591941054458e-06 lb0 = 1.54529351662598e-12 wb0 = 2.30213417558899e-12 pb0 = -1.57695039960758e-18
+ b1 = -3.04989612485908e-09 lb1 = 2.08916359604784e-15 wb1 = 3.11237629687295e-15 pb1 = -2.13196220147648e-21
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0361879334253936+0*(0.009/sqrt(l*w*mult))} lvoff = -4.91249906485148e-08 wvoff = -3.046978156815e-08 pvoff = 3.78501175448116e-14
+ nfactor = {1.43076205861949+0*(0.02/sqrt(l*w*mult))} lnfactor = -8.61735864958842e-08 wnfactor = 3.04139497359176e-07 pnfactor = 9.1898209722022e-14
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -8.03125007569997e-05 lcit = 6.1863611456041e-11 wcit = 6.95845174582576e-11 pcit = -4.76650465363192e-17
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.507529189914283 leta0 = -4.04808253379291e-07 weta0 = -3.63221115474288e-07 peta0 = 3.11899091913197e-13
+ etab = 0.0564211663636824 letab = -4.09331720648957e-08 wetab = -4.68161673670882e-08 petab = 3.15384360115932e-14
+ dsub = 0.880206603104794 ldsub = -5.28411377886793e-07 wdsub = -4.3474741362474e-07 pdsub = 4.07133568902483e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 3.17890110576361 lpclm = -1.42611708945153e-06 wpclm = -1.54724476211258e-06 ppclm = 1.09880325178315e-12
+ pdiblc1 = -2.15888779395002 lpdiblc1 = 1.59465843622959e-06 wpdiblc1 = 2.0845557394419e-06 ppdiblc1 = -1.22866199989679e-12
+ pdiblc2 = -0.0622256668066367 lpdiblc2 = 5.68016672277229e-08 wpdiblc2 = 4.95085960553139e-08 ppdiblc2 = -4.37648893756193e-14
+ pdiblcb = -0.025
+ drout = 9.11531537666202 ldrout = -5.61599460879115e-06 wdrout = -6.69511794621923e-06 pdrout = 4.32704522214906e-12
+ pscbe1 = -396802974.028328 lpscbe1 = 716.170655563672 wpscbe1 = 520.03145411049 ppscbe1 = -0.000551799463722631
+ pscbe2 = 2.71822263184613e-08 lpscbe2 = -1.15565927834355e-14 wpscbe2 = -9.76071644924399e-15 ppscbe2 = 8.90419294733811e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.000887082195626749 lalpha0 = -5.16897396758928e-10 walpha0 = -6.83484335531072e-10 palpha0 = 3.98262207639199e-16
+ alpha1 = -3.081944e-10 walpha1 = 3.145080704784e-16
+ beta0 = 229.663478966301 lbeta0 = -3.09829050710832e-05 wbeta0 = -0.000174641037254829 pbeta0 = 2.38718945965987e-11
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -7.33423919601145e-08 lagidl = 7.14169056985188e-14 wagidl = 5.62359820066937e-14 pagidl = -5.47118470162486e-20
+ bgidl = -304964402.783825 lbgidl = 3038.74059472073 wbgidl = 1027.4156538433 pbgidl = -0.002341307085864
+ cgidl = -3687.96958532273 lcgidl = 0.00185368125366881 wcgidl = 0.00360743824707697 pcgidl = -1.42823545441427e-9
+ egidl = -3.26379626326786 legidl = 7.68552802473515e-07 wegidl = 3.21560045549336e-06 pegidl = -5.92159174566608e-13
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.566951379045799 lkt1 = -3.56026239985612e-08 wkt1 = -6.37662754084442e-08 pkt1 = 2.85990279217913e-14
+ kt2 = -0.019032
+ at = -41306.0615139992 lat = 0.0631055079095819 wat = 0.107718227868675 pat = -9.53300930726383e-8
+ ute = -1.34705075 lute = -9.09325725037485e-8
+ ua1 = 5.524e-10
+ ub1 = -3.5909e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.41e-6
+ sbref = 2.41e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.70 pmos
* DC IV MOS Parameters
+ lmin = 6e-07 lmax = 8.0e-07 wmin = 7.5e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.953287238590066+0*(0.0/sqrt(l*w*mult))} lvth0 = 4.06172509948671e-08 wvth0 = 8.99797170222211e-08 pvth0 = -4.25867648453404e-14
+ k1 = 0.212020778063646 lk1 = 2.86123852192686e-07 wk1 = 2.47717600259682e-07 pk1 = -2.06568038812115e-13
+ k2 = 0.103035847097089 lk2 = -5.52367839692691e-08 wk2 = -5.54489917163869e-08 pk2 = 4.60301349387492e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -140908.778630099 lvsat = 0.109143518874946 wvsat = 0.170723246360216 pvsat = -9.07692562048839e-8
+ ua = -7.01445925326854e-09 lua = 4.35137037725015e-15 wua = 8.9802452531918e-15 pua = -4.72999124348089e-21
+ ub = 1.8402815813418e-17 lub = -9.95142371298983e-24 wub = -1.80719363595758e-23 pub = 1.01406935532887e-29
+ uc = 9.09909918719974e-12 luc = -5.61242060012038e-18 wuc = -9.07591064882698e-18 puc = 4.26273104839137e-24
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0169104816360262 lu0 = -3.28835151756486e-09 wu0 = 1.71744304398526e-09 pu0 = 1.31766795015662e-15
+ a0 = 1.04573163615046 la0 = -5.14211153849152e-08 wa0 = -3.68671473329737e-07 pa0 = 1.30450276407145e-13
+ keta = -0.596203521782092 lketa = 2.96588945700316e-07 wketa = 5.09976984921236e-07 pketa = -2.80402790772956e-13
+ a1 = 0.0
+ a2 = 0.5
+ ags = 5.70122426728559 lags = -2.76100297332191e-06 wags = -5.03371667952024e-06 pags = 2.79462133002893e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.379901736377878+0*(0.009/sqrt(l*w*mult))} lvoff = 1.86317245804922e-07 wvoff = 2.9333030111872e-07 pvoff = -1.83951320095281e-13
+ nfactor = {-4.09506709213075+0*(0.02/sqrt(l*w*mult))} lnfactor = 3.69899175262228e-06 wnfactor = 5.7674844768746e-06 pnfactor = -3.65046578452114e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -2.7368185757e-05 lcit = 2.55970204026162e-11 wcit = 3.81337104104179e-11 pcit = -2.61214009625842e-17
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -0.306661903079854 leta0 = 1.52908574366227e-07 weta0 = 2.92553859637772e-07 peta0 = -1.37303487163689e-13
+ etab = -0.0114247760580253 letab = 5.54095926426199e-09 wetab = -2.6520227701268e-09 petab = 1.28621778339765e-15
+ dsub = -0.146834007263317 ldsub = 1.75106305012311e-07 wdsub = 4.04114410847387e-07 pdsub = -1.67482586551801e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.98276279855881 lpclm = -6.06768329707776e-07 wpclm = -7.16403891869476e-07 ppclm = 5.29681409870976e-13
+ pdiblc1 = 1.11467286848843 lpdiblc1 = -6.47714249737434e-07 wpdiblc1 = -5.36533204703576e-07 ppdiblc1 = 5.66770821398135e-13
+ pdiblc2 = 0.0271736694432785 lpdiblc2 = -4.43643110678779e-09 wpdiblc2 = -2.40710040932812e-08 ppdiblc2 = 6.63676882816762e-15
+ pdiblcb = -0.025
+ drout = 4.24912218893285 ldrout = -2.28267660616261e-06 wdrout = -4.01691669772287e-06 pdrout = 2.49249075793529e-12
+ pscbe1 = 1860384638.62157 lpscbe1 = -829.991573163443 wpscbe1 = -1446.79080263912 ppscbe1 = 0.000795463948039569
+ pscbe2 = -1.1383147601461e-09 lpscbe2 = 7.84283625270517e-15 wpscbe2 = 1.21236140891494e-14 ppscbe2 = -6.08646404980865e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.000416305126641977 lalpha0 = -1.94417458389704e-10 walpha0 = -3.84782790450476e-10 palpha0 = 1.93653142766717e-16
+ alpha1 = -1.05555811514e-09 lalpha1 = 5.11940408052324e-16 walpha1 = 1.07718227868676e-15 palpha1 = -5.22428019251684e-22
+ beta0 = 524.753051998438 lbeta0 = -0.000233117787150232 wbeta0 = -0.000488883768200885 pbeta0 = 2.39126594080992e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -1.41863260421059e-07 lagidl = 1.18353357989923e-13 wagidl = 5.55662806614289e-14 pagidl = -5.42531049432489e-20
+ bgidl = 11827597207.5328 lbgidl = -5272.0034455381 wbgidl = -9651.23430584989 pbgidl = 0.00497351474327603
+ cgidl = -6945.94697927908 lcgidl = 0.00408537947864194 wcgidl = 0.006480247723837 pcgidl = -3.3960955819475e-9
+ egidl = -12.2202832127237 legidl = 6.90370158041599e-06 wegidl = 1.00350022804924e-05 pegidl = -5.26341532768179e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.161452898870202 lkt1 = -3.13367055426447e-07 wkt1 = -4.56739863612253e-07 pkt1 = 2.9778397097346e-13
+ kt2 = -0.019032
+ at = 149805.561514 lat = -0.0678049983064824 wat = -0.107718227868676 pat = 5.22428019251684e-8
+ ute = -1.815901535 lute = 2.30227870967326e-7
+ ua1 = 5.53369990000002e-10 lua1 = -6.64438300050783e-19
+ ub1 = -7.76500946750001e-18 lub1 = 2.85924411469016e-24
+ uc1 = 4.29439976775701e-10 luc1 = -3.68965690891471e-16 wuc1 = -5.49674555339928e-16 puc1 = 3.76524322035074e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.02e-6
+ sbref = 2.01e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.71 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 6e-07 wmin = 7.5e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.02/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.42816446878934+0*(0.0/sqrt(l*w*mult))} lvth0 = -2.14064666744634e-07 wvth0 = -3.60715380786512e-07 pvth0 = 1.75998104116406e-13
+ k1 = 1.4125042238514 lk1 = -2.96104616597147e-07 wk1 = -5.34550586542708e-07 pk1 = 1.72828120446109e-13
+ k2 = -0.10543273735757 lk2 = 4.58694371483178e-08 wk2 = 3.79198373986732e-08 pk2 = 7.46719662090592e-16
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -339935.637967769 lvsat = 0.205670550519419 wvsat = 0.277367723728604 pvsat = -1.42491294506165e-7
+ ua = 1.1796116617539e-08 lua = -4.77166486721217e-15 wua = -1.10707194615981e-14 pua = 4.99462638836861e-21
+ ub = -2.66636704434641e-17 lub = 1.19055967891667e-23 wub = 2.70930849273386e-23 pub = -1.17641159457584e-29
+ uc = 2.11227520703005e-11 luc = -1.14438321301599e-17 wuc = -1.18113460279589e-17 puc = 5.58940353009346e-24
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = -0.00308591797769675 lu0 = 6.40980231309267e-09 wu0 = 1.53437415361241e-08 pu0 = -5.29101868703824e-15
+ a0 = 1.32804257469546 la0 = -1.88340509024551e-07 wa0 = -1.95414274405376e-08 pa0 = -3.88760501988873e-14
+ keta = -0.359550098390452 lketa = 1.81813218622487e-07 wketa = 1.45455556917319e-07 pketa = -1.03611720798197e-13
+ a1 = 0.0
+ a2 = 0.5
+ ags = 9.95408225759512 lags = -4.82361783433208e-06 wags = -7.03850052216094e-06 pags = 3.76693146979045e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {0.62149681335444+0*(0.009/sqrt(l*w*mult))} lvoff = -2.99356043822503e-07 wvoff = -5.85339785337174e-07 pvoff = 2.42199278485395e-13
+ nfactor = {13.5557464269134+0*(0.02/sqrt(l*w*mult))} lnfactor = -4.86156455004654e-06 wnfactor = -1.2334321940736e-05 pnfactor = 5.12881981898791e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 0.000163312773028 lcit = -6.68822912033149e-11 wcit = -1.36809438117752e-10 pcit = 5.87251513578354e-17
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -1.60737052028686 leta0 = 7.83745750168538e-07 weta0 = 1.11419748234508e-06 peta0 = -5.35796535958619e-13
+ etab = 0.120140674511516 letab = -5.82676264347129e-08 wetab = -7.95970118209471e-08 petab = 3.86041527481002e-14
+ dsub = -0.133337343455208 ldsub = 1.68560490548697e-07 wdsub = 3.88389991442807e-07 pdsub = -1.59856321762677e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 5.80914249737145 lpclm = -2.46254335173341e-06 wpclm = -3.00202491153058e-06 ppclm = 1.63819617630151e-12
+ pdiblc1 = -1.01721472019 lpdiblc1 = 3.86240571333659e-07 wpdiblc1 = 2.48882053444533e-06 ppdiblc1 = -9.0051061532039e-13
+ pdiblc2 = 0.0987333941160206 lpdiblc2 = -3.91425397744443e-08 wpdiblc2 = -7.00780178531688e-08 ppdiblc2 = 2.89499404666443e-14
+ pdiblcb = 3.11805606056 lpdiblcb = -1.5243664740913e-06 wpdiblcb = -2.42168069187663e-06 ppdiblcb = 1.17450302715671e-12
+ drout = -6.06868590141123 ldrout = 2.72140872861382e-06 wdrout = 5.44306244123191e-06 pdrout = -2.09555182456208e-12
+ pscbe1 = -7103235374.67175 lpscbe1 = 3517.31931518375 wpscbe1 = 5781.13781088934 ppscbe1 = -0.00271004528987867
+ pscbe2 = 1.58451495433671e-07 lpscbe2 = -6.9557423742245e-14 wpscbe2 = -1.1170401939623e-13 ppscbe2 = 5.39693190524331e-20
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.000242639283311392 lalpha0 = -1.10190392703587e-10 walpha0 = -1.1655357166516e-10 palpha0 = 6.35633128019322e-17
+ alpha1 = 0.0
+ beta0 = 168.446981972935 lbeta0 = -6.03111247182129e-05 wbeta0 = -8.31095598023833e-05 pbeta0 = 4.23281318787605e-11
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 6.9456335031836e-07 lagidl = -2.87309366085641e-13 wagidl = -5.24892158493762e-13 pagidl = 2.27266335754823e-19
+ bgidl = -6344835136.0712 lbgidl = 3541.53537894812 wbgidl = 6100.75615780801 pbgidl = -0.00266612187164573
+ cgidl = 12418.5925977768 lcgidl = -0.00530632539353228 wcgidl = -0.00907061623931866 pcgidl = 4.14599568586318e-9
+ egidl = 18.6704372704376 legidl = -8.07814340031481e-06 wegidl = -1.35796642416696e-05 pegidl = 6.18957986223417e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -2.127281078766 lkt1 = 6.40049782682115e-07 wkt1 = 1.3075523638806e-06 pkt1 = -5.57888937899435e-13
+ kt2 = -0.019032
+ at = 92110.8712112 lat = -0.039823361983076 wat = -0.0484336138375327 pat = 2.34900605431341e-8
+ ute = -3.57029512905663 lute = 1.08109999211682e-06 wute = 1.80173043475621e-06 pute = -8.7383025220459e-13
+ ua1 = 5.52e-10
+ ub1 = -6.90256174897151e-18 lub1 = 2.44096128344244e-24 wub1 = 6.27699635334423e-24 pub1 = -3.04431184639018e-30
+ uc1 = -1.1864799535514e-09 luc1 = 4.14747395717522e-16 wuc1 = 1.09934911067986e-15 puc1 = -4.23243910866191e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 1.81e-6
+ sbref = 1.81e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.72 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 7e-07 wmax = 7.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.911001+0*(0.0/sqrt(l*w*mult))}
+ k1 = 0.57102
+ k2 = 0.0282628
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 180350.0
+ ua = 2.33385448e-9
+ ub = 7.449e-20
+ uc = -3.2639e-11
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.01966047
+ a0 = 0.87668
+ keta = -0.0076977
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.1244
+ b0 = 6.3575e-8
+ b1 = 2.0655e-10
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.10903374+0*(0.009/sqrt(l*w*mult))}
+ nfactor = {1.74899+0*(0.02/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.0800000000000101
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.99495
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00129
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 225600350.0
+ pscbe2 = 1.4994384e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.8978653e-5
+ alpha1 = 0.0
+ beta0 = 37.686511
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 3.08e-8
+ bgidl = 1701900000.0
+ cgidl = 1200.0
+ egidl = 1.0890786
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.566
+ kt2 = -0.019032
+ at = 351440.0
+ ute = -1.4104
+ ua1 = 2.2096e-11
+ ub1 = -2.3998e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.73 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 7e-07 wmax = 7.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.90082738520125+0*(0.0/sqrt(l*w*mult))} lvth0 = -2.02302279405102e-7
+ k1 = 0.5619325432625 lk1 = 1.80704031787894e-7
+ k2 = 0.0309775045589796 lk2 = -5.39818865817867e-8
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 246185.7657525 lvsat = -1.30914387280963
+ ua = 2.38881257975021e-09 lua = -1.09284153874223e-15
+ ub = -9.53776338333291e-21 lub = 1.67089165473876e-24 pub = 1.40129846432482e-45
+ uc = -2.4445450689826e-11 luc = -1.62928687065067e-16
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.02024593087875 lu0 = -1.16418866466391e-8
+ a0 = 0.857053117262389 la0 = 3.90280465103088e-7
+ keta = -0.00737954045175002 lketa = -6.3266010261535e-9
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.1232871118057 lags = 2.21297761792142e-8
+ b0 = 1.05349046427083e-07 lb0 = -8.3067670433232e-13
+ b1 = 3.42270476437501e-10 lb1 = -2.69880099535731e-15
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.109923174006829+0*(0.009/sqrt(l*w*mult))} lvoff = 1.76863907786298e-8
+ nfactor = {1.81308843852084+0*(0.02/sqrt(l*w*mult))} lnfactor = -1.27459712949456e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.32854145833333e-05 lcit = -6.53304525625104e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.0800000000000101
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.59382769055469 lpclm = -1.19086798822915e-5
+ pdiblc1 = 0.39
+ pdiblc2 = -0.000121457866722241 lpdiblc2 = 2.80668326224826e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 226180383.373859 lpscbe1 = -11.5339607389978
+ pscbe2 = 1.49915329172246e-08 lpscbe2 = 5.66937667336574e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -1.07635402550049e-05 lalpha0 = 5.91423364164808e-10
+ alpha1 = 0.0
+ beta0 = 36.7974994974862 lbeta0 = 1.76779892824275e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 3.78964955000001e-08 lagidl = -1.41113777535023e-13
+ bgidl = 1821160549.375 lbgidl = -2371.49542801909
+ cgidl = 1068.58341666667 lcgidl = 0.00261321810250043
+ egidl = 0.805970088606919 legidl = 5.6296113335089e-6
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.572570829166667 lkt1 = 1.30660905125007e-7
+ kt2 = -0.019032
+ at = 483086.562354168 lat = -2.61779123417979
+ ute = -1.31466301904167 lute = -1.90372938767156e-6
+ ua1 = 2.2096e-11
+ ub1 = -1.95502057370835e-18 lub1 = -8.84443666791263e-24
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.74 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 7e-07 wmax = 7.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.941521844396252+0*(0.0/sqrt(l*w*mult))} lvth0 = 1.18573327875207e-7
+ k1 = 0.598282370212502 lk1 = -1.05914171963714e-7
+ k2 = 0.0201186863230615 lk2 = 3.16398409143385e-8
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -17157.2972574998 lvsat = 0.767314862308899 pvsat = -8.470329472543e-22
+ ua = 2.1689801807494e-09 lua = 6.40535828217084e-16
+ ub = 3.2657329015e-19 lub = -9.793423218163e-25
+ uc = -5.72196479305226e-11 luc = 9.54956943068406e-17
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0179040873637502 lu0 = 6.82353775991796e-9
+ a0 = 0.935560648212853 la0 = -2.28751023903696e-7
+ keta = -0.00865217864475001 lketa = 3.70814476246048e-9
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.127738664582901 lags = -1.29706952112439e-8
+ b0 = -6.174713928125e-08 lb0 = 4.86875884496959e-13
+ b1 = -2.006114293125e-10 lb1 = 1.58182011707191e-15
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.106365437979512+0*(0.009/sqrt(l*w*mult))} lvoff = -1.03663400080826e-8
+ nfactor = {1.5566946844375+0*(0.02/sqrt(l*w*mult))} lnfactor = 7.47066339483736e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.43756250000016e-07 lcit = 3.82914576875313e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.0800000000000101
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.801683071664061 lpclm = 6.97991050024954e-06 wpclm = 4.2351647362715e-22 ppclm = 1.61558713389263e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00552437360016675 lpdiblc2 = -1.64505202647799e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 223860249.878426 lpscbe1 = 6.76028027181746
+ pscbe2 = 1.50029372483263e-08 lpscbe2 = -3.3229326980971e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.000108205232765015 lalpha0 = -3.46644816254184e-10 palpha0 = 7.88860905221012e-31
+ alpha1 = 0.0
+ beta0 = 40.3535455075414 lbeta0 = -1.03614157266245e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 9.51051350000005e-09 lagidl = 8.27095486050672e-14
+ bgidl = 1344118351.87502 lbgidl = 1389.97991405736
+ cgidl = 1594.24975 lcgidl = -0.00153165830750124
+ egidl = 1.93840413417926 legidl = -3.29962545365871e-6
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.546287512500001 lkt1 = -7.65829153750579e-8
+ kt2 = -0.019032
+ at = -43499.6870625 lat = 1.53433870953938
+ ute = -1.697610942875 lute = 1.11581307701467e-6
+ ua1 = 2.2096e-11
+ ub1 = -3.73413827887501e-18 lub1 = 5.183897541738e-24
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.75 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 7e-07 wmax = 7.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.93885745611+0*(0.0/sqrt(l*w*mult))} lvth0 = 1.08222192705071e-7
+ k1 = 0.58155712205 lk1 = -4.09366664786385e-8
+ k2 = 0.0220218228343599 lk2 = 2.42461650836256e-8
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 314326.019625001 lvsat = -0.520496166363026 pvsat = 8.470329472543e-22
+ ua = 2.61942847040729e-09 lua = -1.10945352486243e-15
+ ub = 3.84703627149999e-19 lub = -1.20517839040961e-24 wub = -3.67341984631965e-40 pub = -7.00649232162409e-46
+ uc = -6.07650070962588e-11 luc = 1.0926939693893e-16
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0216706946428249 lu0 = -7.80971268625172e-9
+ a0 = 1.00612260665 la0 = -5.02883879622213e-7
+ keta = 0.02009777652175 lketa = -1.07985287309616e-07 pketa = -5.04870979341448e-29
+ a1 = 0.0
+ a2 = 0.5
+ ags = -0.165909842420324 lags = 1.12785228625375e-6
+ b0 = 3.43010276499998e-08 lb0 = 1.13729236209888e-13
+ b1 = 3.4088605367e-10 lb1 = -5.2189489682768e-16
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.140418550485945+0*(0.009/sqrt(l*w*mult))} lvoff = 1.21929831813844e-7
+ nfactor = {1.581762668575+0*(0.02/sqrt(l*w*mult))} lnfactor = 6.49677346449464e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.0988499500000101 leta0 = -7.32319615002507e-8
+ etab = -0.135974825 letab = 2.56311865250875e-7
+ dsub = 0.790011133214275 ldsub = -8.93592102481797e-07 wdsub = -1.6940658945086e-21
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.829249703024498 lpclm = 6.43744825248333e-7
+ pdiblc1 = 0.242386211199548 lpdiblc1 = 5.73478831420806e-7
+ pdiblc2 = 0.0005919348911365 lpdiblc2 = 2.71197945760915e-9
+ pdiblcb = -0.025
+ drout = 0.686444022578826 ldrout = -4.91234395498629e-7
+ pscbe1 = 176085112.8405 lpscbe1 = 192.366448788471
+ pscbe2 = 1.54471758214575e-08 lpscbe2 = -1.75909396240323e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.68658917561175e-05 lalpha0 = -6.94918331313226e-11
+ alpha1 = -9.42497500000001e-11 lalpha1 = 3.6615980750125e-16
+ beta0 = 70.3784609012225 lbeta0 = -0.0001270080619065
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 5.97293952639999e-08 lagidl = -1.12390555953664e-13
+ bgidl = 2336577816.5 lbgidl = -2465.72014371341
+ cgidl = 757.026174999992 lcgidl = 0.00172095109525587
+ egidl = 1.25816693043865 legidl = -6.56907318312498e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.488715204999995 lkt1 = -3.00251042151023e-7
+ kt2 = -0.019032
+ at = 649872.408399999 lat = -1.15940841447196
+ ute = -1.3732655985 lute = -1.44266964155498e-7
+ ua1 = -4.77714194239999e-10 lua1 = 1.94176010557143e-15 pua1 = 1.88079096131566e-37
+ ub1 = -1.27719122775e-18 lub1 = -4.36132946714737e-24
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.76 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 7e-07 wmax = 7.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.90159456616+0*(0.0/sqrt(l*w*mult))} lvth0 = 3.79818314637668e-8
+ k1 = 0.55984
+ k2 = 0.0353628837975001 lk2 = -9.01668126588628e-10
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 10474.8766399999 lvsat = 0.0522617189079835
+ ua = 2.031112101561e-09 lua = -4.80111168975445e-19
+ ub = -2.8312028915e-19 lub = 5.36663526963041e-26
+ uc = -2.7970035e-12
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0177626546720001 lu0 = -4.43076881446636e-10
+ a0 = 0.73934
+ keta = -0.041230772165 lketa = 7.61872032216419e-9
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.43242187
+ b0 = 3.1990628925e-08 lb0 = 1.1808432625452e-13
+ b1 = -7.72466718899999e-11 lb1 = 2.66283200189291e-16
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.075734118+0*(0.009/sqrt(l*w*mult))}
+ nfactor = {1.98263488240001+0*(0.02/sqrt(l*w*mult))} lnfactor = -1.05964772249584e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.0811416455550104 leta0 = -3.98518961629476e-8
+ etab = 0.00384149779649999 letab = -7.24120413891353e-9
+ dsub = 0.31595571
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.1707598
+ pdiblc1 = 0.54661982
+ pdiblc2 = 0.0020306546
+ pdiblcb = -0.025
+ drout = 0.42584153
+ pscbe1 = 278136550.0
+ pscbe2 = 1.4513967e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 3.0
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.056e-10
+ bgidl = 1028500000.0
+ cgidl = 2268.2035203 lcgidl = -0.0011276106447479
+ egidl = 0.90967406
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.648
+ kt2 = -0.019032
+ at = 39047.976 lat = -0.00800741352011991
+ ute = -1.4498
+ ua1 = 5.524e-10
+ ub1 = -3.5909e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.81e-6
+ sbref = 2.81e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.77 pmos
* DC IV MOS Parameters
+ lmin = 8.0e-07 lmax = 1e-06 wmin = 7e-07 wmax = 7.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.861341630549994+0*(0.0/sqrt(l*w*mult))} lvth0 = 2.35818471359657e-9
+ k1 = 0.55984
+ k2 = 0.0230344340525002 lk2 = 1.00089482554878e-8
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 74688.7523299996 lvsat = -0.00456724000828856
+ ua = 2.02846050039498e-09 lua = 1.86654260492757e-18
+ ub = 2.69962905500005e-19 lub = -4.35809509152973e-25
+ uc = -2.7970035e-12
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0187224093399998 lu0 = -1.29245496385334e-9
+ a0 = 0.73934
+ keta = -0.032622
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.43242187
+ b0 = 7.31979364499999e-07 lb0 = -5.01402204785677e-13
+ b1 = 9.89601408999999e-10 lb1 = -6.77872017157955e-16
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.075734118+0*(0.009/sqrt(l*w*mult))}
+ nfactor = {1.82549927299999+0*(0.02/sqrt(l*w*mult))} lnfactor = 3.30994563913558e-8
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.0361110000000101
+ etab = -0.0043407
+ dsub = 0.31595571
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.1707598
+ pdiblc1 = 0.54661982
+ pdiblc2 = 0.0020306546
+ pdiblcb = -0.025
+ drout = 0.42584153
+ pscbe1 = 278136550.0
+ pscbe2 = 1.4513967e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 3.0
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -3.5471664e-10 lagidl = 4.07377924816799e-16
+ bgidl = 1028500000.0
+ cgidl = 994.06
+ egidl = 0.90967406
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.649712487500004 lkt1 = 1.51554287506185e-9
+ kt2 = -0.019032
+ at = 98499.4999999998 lat = -0.0606217150024999
+ ute = -1.34705074999998 lute = -9.09325725037519e-8
+ ua1 = 5.524e-10
+ ub1 = -3.5909e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.41e-6
+ sbref = 2.41e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.78 pmos
* DC IV MOS Parameters
+ lmin = 6e-07 lmax = 8.0e-07 wmin = 7e-07 wmax = 7.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.014/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.836504173067496+0*(0.0/sqrt(l*w*mult))} lvth0 = -1.46553494746287e-8
+ k1 = 0.533529021250001 lk1 = 1.80228888888591e-8
+ k2 = 0.0310695924001998 lk2 = 4.50490496310518e-9
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 80669.8695999999 lvsat = -0.00866427543265202
+ ua = 4.64084045781224e-09 lua = -1.78760066632611e-15
+ ub = -5.05242718850001e-18 lub = 3.21000109328656e-24 wub = 5.87747175411144e-39 pub = 1.40129846432482e-45
+ uc = -2.68036292999249e-12 luc = -7.98982072522827e-20
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.019139520248 lu0 = -1.57817385027881e-9
+ a0 = 0.567239524250006 la0 = 1.17887965386369e-7
+ keta = 0.0656864865000002 lketa = -6.73408217100675e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = -0.831946587889249 lags = 8.66086071811846e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {0.000806415514200687+0*(0.009/sqrt(l*w*mult))} lvoff = -5.24298827545597e-8
+ nfactor = {3.3904478645+0*(0.02/sqrt(l*w*mult))} lnfactor = -1.03888250404318e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 2.21248750000001e-05 lcit = -8.30547875062503e-12 wcit = -5.16987882845642e-26
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.0730385193000101 leta0 = -2.52951660829035e-8
+ etab = -0.0148667889825 letab = 7.2103183225676e-9
+ dsub = 0.377658859378499 ldsub = -4.2266348808525e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.05295499949499 lpclm = 8.06956993219213e-8
+ pdiblc1 = 0.418316017483253 lpdiblc1 = 8.78874632049621e-8
+ pdiblc2 = -0.00406765628266752 lpdiblc2 = 4.17731246307284e-9
+ pdiblcb = -0.025
+ drout = -0.964362154355499 ldrout = 9.52282572765097e-7
+ pscbe1 = -17379269.6637516 lpscbe1 = 202.426858890571
+ pscbe2 = 1.4596707147e-08 lpscbe2 = -5.66765869943222e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -8.30975756141003e-05 lalpha0 = 5.69214923072805e-11 walpha0 = -4.8778425213436e-26 palpha0 = -3.6055891202998e-32
+ alpha1 = 3.424975e-10 lalpha1 = -1.661095750125e-16
+ beta0 = -109.760447534175 lbeta0 = 7.72403427586724e-05 wbeta0 = 2.71050543121376e-20 pbeta0 = 5.16987882845642e-26
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -6.97447785e-08 lagidl = 4.79392233486075e-14 wagidl = 1.57772181044202e-30 pagidl = -2.25694915357879e-36
+ bgidl = -698567194.999992 lbgidl = 1183.03239323903
+ cgidl = 1464.6506485 lcgidl = -0.000322352241269259
+ egidl = 0.803966780776996 legidl = 7.24089577313559e-8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.754247399500002 lkt1 = 7.31214349205069e-8
+ kt2 = -0.019032
+ at = 10000.0
+ ute = -1.81590153499999 lute = 2.30227870967324e-7
+ ua1 = 5.53369989999999e-10 lua1 = -6.64438300050783e-19
+ ub1 = -7.76500946749999e-18 lub1 = 2.85924411469015e-24
+ uc1 = -2.83972798199999e-10 luc1 = 1.19718492903009e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.02e-6
+ sbref = 2.01e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.79 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 6e-07 wmin = 7e-07 wmax = 7.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.896330510464999+0*(0.0/sqrt(l*w*mult))} lvth0 = 1.43601250314735e-8
+ k1 = 0.718720577499994 lk1 = -7.17940899346127e-8
+ k2 = -0.0562172585576 lk2 = 4.68385912433833e-8
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 20054.9702049997 lvsat = 0.020733647699426
+ ua = -2.57237218251451e-09 lua = 1.71077139816917e-15
+ ub = 8.49995995e-18 lub = -3.36283890695025e-24
+ uc = 5.79301729516001e-12 luc = -4.18944524955012e-18
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0168284497540001 lu0 = -4.57316216041203e-10
+ a0 = 1.3026801055 la0 = -2.38797039316976e-7
+ keta = -0.1707659324 lketa = 4.7337419194338e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.818938306684998 lags = 6.5415152367809e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.138205225796401+0*(0.009/sqrt(l*w*mult))} lvoff = 1.49900682228749e-8
+ nfactor = {-2.45274943250001+0*(0.02/sqrt(l*w*mult))} lnfactor = 1.79503896901534e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -1.42497500000001e-05 lcit = 9.33603250125e-12
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -0.161273534299991 leta0 = 8.83450083528289e-08 peta0 = 1.0097419586829e-28
+ etab = 0.016833136385 letab = -8.1639869810431e-9
+ dsub = 0.370747080457498 ldsub = -3.89141705907336e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.91286805302001 lpclm = -3.36357832072436e-7
+ pdiblc1 = 2.2129809413085 lpdiblc1 = -7.82516051525667e-7
+ pdiblc2 = 0.00778038802224501 lpdiblc2 = -1.56892978458824e-9
+ pdiblcb = -0.025
+ drout = 0.995767497134494 ldrout = 1.62949244070272e-9
+ pscbe1 = 400000000.0
+ pscbe2 = 1.34728463781e-08 lpscbe2 = 4.88390266618356e-16
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 9.13664870955504e-05 lalpha0 = -2.76927057865862e-11
+ alpha1 = 0.0
+ beta0 = 60.5805706398501 lbeta0 = -5.37419935063913e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.33152049999999e-08 lagidl = 7.65554665102504e-15
+ bgidl = 1573227175.0 lbgidl = 81.2234827608772
+ cgidl = 646.002 lcgidl = 7.46882600100029e-5
+ egidl = 1.04563391038999 legidl = -4.47983917952942e-8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.430232249999996 lkt1 = -8.40242925112479e-8
+ kt2 = -0.019032
+ at = 29249.75 lat = -0.00933603250124998
+ ute = -1.23186141999999 lute = -5.30286646070998e-8
+ ua1 = 5.52e-10
+ ub1 = 1.24423955999998e-18 lub1 = -1.5101966174022e-24
+ uc1 = 2.403455964e-10 luc1 = -1.34573306886018e-16 puc1 = 9.4039548065783e-38
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 1.81e-6
+ sbref = 1.81e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.80 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 4.2e-07 wmax = 7.0e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.85055751108+0*(0.0/sqrt(l*w*mult))} wvth0 = -4.35486875580151e-8
+ k1 = 0.521009107357143 wk1 = 3.60321479966816e-8
+ k2 = 0.0411922785828286 wk2 = -9.31550830622783e-9
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 422036.802378571 wvsat = -0.174131957498527
+ ua = 3.514423473386e-09 wua = -8.50583431768705e-16
+ ub = -1.29257403264286e-18 wub = 9.84950496622721e-25
+ uc = -1.83661162022214e-11 wuc = -1.02834129559263e-17
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0200931216418571 wu0 = -3.11719450835086e-10
+ a0 = 0.833150544214286 wa0 = 3.13623634812261e-8
+ keta = -0.0131943360142857 wketa = 3.96024929538866e-9
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.1504929590605 wags = -1.87996117016634e-8
+ b0 = 1.53287997037857e-07 wb0 = -6.46369583838175e-14
+ b1 = -1.61770907953571e-08 wb1 = 1.18041838220837e-14
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0883533942492857+0*(0.009/sqrt(l*w*mult))} wvoff = -1.48998995885491e-8
+ nfactor = {1.77257173264286+0*(0.02/sqrt(l*w*mult))} wnfactor = -1.6990308224922e-8
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 2.55871059043665e-05 wcit = -1.12302915846134e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.0800000000000101
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.42876142683036 wpclm = -1.0330410596713e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00129
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 226544799.178928 wpscbe1 = -0.680462411129554
+ pscbe2 = 1.49855491093714e-08 wpscbe2 = 6.36541500941602e-18
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 4.88350347741357e-05 walpha0 = -2.15111050789199e-11
+ alpha1 = -1.57316428571429e-10 walpha1 = 1.13344284355714e-16
+ beta0 = 92.2540913012357 wbeta0 = -3.93151776609161e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 6.35218171428571e-08 wagidl = -2.35756111459886e-14
+ bgidl = 2418633648.57143 wbgidl = -516.396559524634
+ cgidl = 885.367142857143 wcgidl = 0.000226688568711428
+ egidl = -0.343950413572857 wegidl = 1.03247734187305e-6
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.582156397214286 wkt1 = 1.16404580033318e-8
+ kt2 = -0.019032
+ at = 830688.768 wat = -0.345292027861248
+ ute = -1.35628314857143 wute = -3.89904338183658e-8
+ ua1 = -1.05467831965714e-09 wua1 = 7.75800822472496e-16
+ ub1 = -1.22747797428572e-18 wub1 = -8.44641607018783e-25
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.81 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 4.2e-07 wmax = 7.0e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.81953769441994+0*(0.0/sqrt(l*w*mult))} lvth0 = -6.1682889918621e-07 wvth0 = -5.85680841522629e-08 pvth0 = 2.98660626179634e-13
+ k1 = 0.448545541800263 lk1 = 1.44093763878073e-06 wk1 = 8.16937471355211e-08 pk1 = -9.07980670567835e-13
+ k2 = 0.0614924020252604 lk2 = -4.03667853152141e-07 wk2 = -2.19855564158908e-08 pk2 = 2.51943843310408e-13
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 646680.837157823 lvsat = -4.46704550836525 wvsat = -0.288551092016536 pvsat = 2.27522391779493e-6
+ ua = 4.30585384311616e-09 lua = -1.57375889449324e-14 wua = -1.38120139167749e-15 pua = 1.05513354796963e-20
+ ub = -2.19162527448937e-18 lub = 1.78776294488617e-23 wub = 1.57216350252674e-24 pub = -1.16767276863364e-29
+ uc = 1.32255337903839e-11 luc = -6.28199802144707e-16 wuc = -2.71414169242084e-17 puc = 3.3522132461927e-22
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0234626037053875 lu0 = -6.70021339858907e-08 wu0 = -2.31756773817274e-09 pu0 = 3.98862831644678e-14
+ a0 = 0.757476770677838 la0 = 1.50477260840339e-06 wa0 = 7.17433636453126e-08 pa0 = -8.02975986357855e-13
+ keta = -0.0133567433065206 lketa = 3.22946819405465e-09 wketa = 4.30649097602226e-09 pketa = -6.88501408819089e-15
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.159306282843203 lags = -1.75252899352433e-07 wags = -2.59513084641265e-08 pags = 1.42211454363095e-13
+ b0 = 2.92438695570863e-07 lb0 = -2.76701094457533e-12 wb0 = -1.34795472953005e-13 pb0 = 1.39510171141573e-18
+ b1 = -1.72264549699713e-08 lb1 = 2.0866601365382e-14 wb1 = 1.26580207219813e-14 pb1 = -1.69785424852796e-20
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0957873857533789+0*(0.009/sqrt(l*w*mult))} lvoff = 1.47824883888936e-07 wvoff = -1.01846375355753e-08 pvoff = -9.37629623470737e-14
+ nfactor = {1.89708989976413+0*(0.02/sqrt(l*w*mult))} lnfactor = -2.47604313061562e-06 wnfactor = -6.05218768053359e-08 pnfactor = 8.65625023563694e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 3.65302930546007e-05 lcit = -2.17605221766472e-10 wcit = -1.67476095102495e-11 pcit = 1.09711839364685e-16
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.0800000000000101
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 3.96977185325189 lpclm = -3.064298462434e-05 wpclm = -1.71183450600505e-06 ppclm = 1.34978042863795e-11
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00215704204427687 lpdiblc2 = -1.72411267152352e-08 wpdiblc2 = -1.64162728687611e-09 ppdiblc2 = 3.2643750391395e-14
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 228037320.341063 lpscbe1 = -29.6787758464416 wpscbe1 = -1.33789708775356 ppscbe1 = 1.30730852574952e-5
+ pscbe2 = 1.49782128049981e-08 lpscbe2 = 1.45882375781908e-16 wpscbe2 = 9.59695437760349e-18 ppscbe2 = -6.42591441786614e-23
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -2.76965146884555e-05 lalpha0 = 1.52182947840588e-09 walpha0 = 1.2199971017659e-11 palpha0 = -6.70344579625092e-16
+ alpha1 = -1.57316428571429e-10 walpha1 = 1.13344284355714e-16
+ beta0 = 89.9665186533781 lbeta0 = 4.54883706647847e-05 wbeta0 = -3.83075339355519e-05 pbeta0 = -2.00369904406483e-11
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.43804228552368e-07 lagidl = -1.59641534946606e-12 wagidl = -7.63050389559683e-14 pagidl = 1.04852440835431e-18
+ bgidl = 2781020291.47633 lbgidl = -7206.05658223072 wbgidl = -691.565506147618 pbgidl = 0.0034832336277533
+ cgidl = 635.075131139717 lcgidl = 0.00497705540154095 wcgidl = 0.000312336650606169 pcgidl = -1.70311168023651e-9
+ egidl = -1.07243512407128 legidl = 1.44859148258375e-05 wegidl = 1.35336465806166e-06 pegidl = -6.38084267797385e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.589006325212811 lkt1 = 1.36210784001029e-07 wkt1 = 1.18415448043022e-08 pkt1 = -3.99861003185864e-15
+ kt2 = -0.019032
+ at = 1277241.50864051 lat = -8.87969901487291 wat = -0.572177520630065 pat = 4.51161688928046e-6
+ ute = -1.22498690903559 lute = -2.6108250666889e-06 wute = -6.46103817938359e-08 pute = 5.09452537392487e-13
+ ua1 = -1.76220833020922e-09 lua1 = 1.40692307221781e-14 wua1 = 1.28556628965512e-15 pua1 = -1.01366837660992e-20
+ ub1 = -1.23857720651302e-20 lub1 = -2.41621023656953e-23 wub1 = -1.3996411776967e-24 pub1 = 1.10361636879326e-29
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.82 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 4.2e-07 wmax = 7.0e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.936723534720365+0*(0.0/sqrt(l*w*mult))} lvth0 = 3.0718086565344e-07 wvth0 = -3.45711494513982e-09 pvth0 = -1.35889090463684e-13
+ k1 = 0.719545100367592 lk1 = -6.95892525524866e-07 wk1 = -8.73680993985216e-08 pk1 = 4.25071144043863e-13
+ k2 = -0.0205469136745409 lk2 = 2.43211740944215e-07 wk2 = 2.92989954798724e-08 pk2 = -1.52434591964925e-13
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -109016.680081704 lvsat = 1.49162563658083 wvsat = 0.0661833992934794 pvsat = -5.21855772512088e-7
+ ua = 1.94952735794828e-09 lua = 2.84203360898389e-15 wua = 1.58112686488685e-16 pua = -1.58614833007355e-21
+ ub = 7.56733526669673e-19 lub = -5.37016495648336e-24 wub = -3.09924428169113e-25 pub = 3.16352623676073e-30
+ uc = -9.13600880648434e-11 luc = 1.96457303255651e-16 wuc = 2.45977091506163e-17 puc = -7.27414257850927e-23
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0137097017712306 lu0 = 9.8994490004265e-09 wu0 = 3.02199609801191e-09 pu0 = -2.21615098602894e-15
+ a0 = 0.916011306449316 la0 = 2.54728586517965e-07 wa0 = 1.4085027049842e-08 pa0 = -3.48340290594251e-13
+ keta = -0.0140151783031798 lketa = 8.42122485053737e-09 wketa = 3.86396617190346e-09 pketa = -3.39570822033815e-15
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.134787028567623 lags = 1.8081298014242e-08 wags = -5.07824757389736e-09 pags = -2.23725263910572e-14
+ b0 = -2.02004541042988e-07 lb0 = 1.1316715039087e-12 wb0 = 1.01053494365707e-13 pb0 = -4.64566216647488e-19
+ b1 = -2.28899777271175e-08 lb1 = 6.55234499878661e-14 wb1 = 1.63473707664404e-14 pb1 = -4.6069049139089e-20
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.104486717868967+0*(0.009/sqrt(l*w*mult))} lvoff = 2.16419074123686e-07 wvoff = -1.35359153756671e-09 pvoff = -1.63395715886142e-13
+ nfactor = {0.633445977718379+0*(0.02/sqrt(l*w*mult))} lnfactor = 7.48778287649549e-06 wnfactor = 6.65187767709232e-07 pnfactor = -4.85659189488546e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 2.56832349174111e-07 lcit = 6.84108345285132e-11 wcit = -8.14697463895569e-14 pcit = -2.17005893426517e-17
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.0800000000000101
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.341512626455649 lpclm = 3.35147194173155e-06 wpclm = -3.31546363386428e-07 ppclm = 2.61423918327238e-12
+ pdiblc1 = 0.39
+ pdiblc2 = -0.0013111261328306 lpdiblc2 = 1.01053620204162e-08 wpdiblc2 = 4.92488186062833e-09 ppdiblc2 = -1.91331414041317e-14
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 222069435.917263 lpscbe1 = 17.3779629958017 wpscbe1 = 1.29025638762175 ppscbe1 = -7.64989175507168e-6
+ pscbe2 = 1.50075748297637e-08 lpscbe2 = -8.56370426845939e-17 wpscbe2 = -3.34131249953372e-18 ppscbe2 = 3.77590254562118e-23
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.000312136316347792 lalpha0 = -1.15775069515078e-09 walpha0 = -1.46929490686221e-10 palpha0 = 5.84390430262694e-16
+ alpha1 = -3.10109813175893e-10 lalpha1 = 1.20477507363928e-15 walpha1 = 2.23429778855846e-16 palpha1 = -8.68023573706068e-22
+ beta0 = 151.010964609404 lbeta0 = -0.00043584678047625 wbeta0 = -7.97271212590247e-05 pbeta0 = 3.06556248506998e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -9.52753695530776e-08 lagidl = 2.88726086197384e-13 wagidl = 7.54967617373797e-14 pagidl = -1.48432031103738e-19
+ bgidl = 1850571825.60455 lbgidl = 130.524918925916 wbgidl = -364.89263747351 pbgidl = 0.000907419691622292
+ cgidl = 1330.65640880049 lcgidl = -0.000507599494907866 wcgidl = 0.000189915312027469 pcgidl = -7.37820037650158e-10
+ egidl = 0.816512063517655 legidl = -4.08424303565282e-07 wegidl = 8.08307530422691e-07 pegidl = -2.08306995182622e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.577298493817589 lkt1 = 4.3894591988867e-08 wkt1 = 2.23429778855847e-08 pkt1 = -8.68023573706063e-14
+ kt2 = -0.019032
+ at = -244866.088632723 lat = 3.12211177908858 wat = 0.145081673201724 pat = -1.14396826778723e-6
+ ute = -1.74650482594843 lute = 1.50134110057922e-06 wute = 3.5227358240042e-08 pute = -2.7776754358594e-13
+ ua1 = 2.2096e-11
+ ub1 = -3.734138278875e-18 lub1 = 5.18389754173799e-24
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.83 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 4.2e-07 wmax = 7.0e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.9208338984315+0*(0.0/sqrt(l*w*mult))} lvth0 = 2.4544970811938e-07 wvth0 = -1.29857209775518e-08 pvth0 = -9.88705036707964e-14
+ k1 = 0.568899787909994 lk1 = -1.10636239853663e-07 wk1 = 9.11943204519601e-09 pk1 = 5.02175668226762e-14
+ k2 = 0.0242987526131503 lk2 = 6.89865516448657e-08 wk2 = -1.64049602860152e-09 pk2 = -3.22348221519617e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 635417.255874051 lvsat = -1.4004964824376 wvsat = -0.231341740440134 pvsat = 6.34027907727302e-7
+ ua = 3.18395901901341e-09 lua = -1.95372722209581e-15 wua = -4.06736356843019e-16 pua = 6.0828737902491e-22
+ ub = 6.18101715930773e-19 lub = -4.83158106492179e-24 wub = -1.68160055393304e-25 pub = 2.61277235734858e-30
+ uc = -8.95016427734455e-11 luc = 1.89237252590797e-16 wuc = 2.07043436925136e-17 puc = -5.7615720447191e-23
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0220201351733954 lu0 = -2.23865432148165e-08 wu0 = -2.51767010108541e-10 pu0 = 1.05024023202034e-14
+ a0 = 1.41844492549922 la0 = -1.69722351132282e-06 wa0 = -2.970724582184e-07 pa0 = 8.60504983885441e-13
+ keta = 0.0538326294590925 lketa = -2.55167169066852e-07 wketa = -2.43054892534142e-08 pketa = 1.06042485259744e-13
+ a1 = 0.0
+ a2 = 0.5
+ ags = -0.629575455390714 lags = 2.98762572637996e-06 wags = 3.34064582826584e-07 pags = -1.33994072678278e-12
+ b0 = 4.27513404601529e-10 lb0 = 3.45223984540089e-13 wb0 = 2.44053927846102e-14 pb0 = -1.66788725245433e-19
+ b1 = -2.43912399037874e-09 lb1 = -1.39280145250954e-14 wb1 = 2.0029583165965e-15 pb1 = 9.65892150649209e-21
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.125469121995106+0*(0.009/sqrt(l*w*mult))} lvoff = 2.97935609241715e-07 wvoff = -1.07708539356507e-08 pvoff = -1.26809698555897e-13
+ nfactor = {2.20047107492872+0*(0.02/sqrt(l*w*mult))} lnfactor = 1.39989820895881e-06 wnfactor = -4.45770744860166e-07 pnfactor = -5.40523628345903e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.78658214285714e-05 wcit = -5.66721421778571e-12
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.73641241474126 leta0 = -2.55015894920768e-06 weta0 = -4.59354829971564e-07 peta0 = 1.78459121766538e-12
+ etab = -1.70245097383519 letab = 6.34206387109483e-06 wetab = 1.12862413456967e-06 petab = -4.38469911968249e-12
+ dsub = 0.707045411391143 ldsub = -5.71270688027536e-07 wdsub = 5.97756410534608e-08 pdsub = -2.3222806661449e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.949825386783475 lpclm = -1.66536978301239e-06 wpclm = -8.68730920887701e-08 ppclm = 1.66368474764734e-12
+ pdiblc1 = 0.296929754193334 lpdiblc1 = 3.61577439607668e-07 wpdiblc1 = -3.92978591174196e-08 ppdiblc1 = 1.5267198618188e-13
+ pdiblc2 = -0.000506236207230813 lpdiblc2 = 6.97836868391068e-09 wpdiblc2 = 7.91216901978272e-10 ppdiblc2 = -3.07387370810108e-15
+ pdiblcb = -0.025
+ drout = 0.515103721387208 ldrout = 1.74421817929305e-07 wdrout = 1.23448288244344e-07 pdrout = -4.79595982587833e-13
+ pscbe1 = 199716558.290353 lpscbe1 = 104.218780811957 wpscbe1 = -17.0261256063831 ppscbe1 = 6.35091607097273e-5
+ pscbe2 = 1.5767618708247e-08 lpscbe2 = -3.0384037103729e-15 wpscbe2 = -2.30874613731433e-16 ppscbe2 = 9.21724763075622e-22
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.60027087857186e-05 lalpha0 = -8.49730104401625e-11 walpha0 = 6.21911245610821e-13 palpha0 = 1.11539715145367e-17
+ alpha1 = -2.425200906375e-10 lalpha1 = 9.42189339526234e-16 walpha1 = 1.0682670464455e-16 palpha1 = -4.15021213410553e-22
+ beta0 = 120.43542123515 lbeta0 = -0.000317060947344991 wbeta0 = -3.60653391231502e-05 pbeta0 = 1.36930443218036e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 6.07482283918743e-08 lagidl = -3.17424811700765e-13 wagidl = -7.34055004969681e-16 pagidl = 1.47724310786206e-19
+ bgidl = 3491964205.55071 lbgidl = -6246.27627020302 wbgidl = -832.439717901591 pbgidl = 0.00272383776134999
+ cgidl = -11.0141895022498 lcgidl = 0.0047047840711453 wcgidl = 0.000553362330058768 pcgidl = -2.14980988546666e-9
+ egidl = 1.36432580991769 legidl = -2.53667796926068e-06 wegidl = -7.64859864403345e-08 pegidl = 1.35434843721905e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.3997530006175 lkt1 = -6.45868761366015e-07 wkt1 = -6.409602278673e-08 pkt1 = 2.49012728046332e-13
+ kt2 = -0.019032
+ at = 1273824.5597716 lat = -2.77799379650896 wat = -0.449548789733117 pat = 1.16616810756231e-6
+ ute = -1.12750403239692 lute = -9.0347388736442e-07 wute = -1.77067767715345e-07 pute = 5.46997959275108e-13
+ ua1 = -4.7771419424e-10 lua1 = 1.94176010557143e-15 wua1 = -1.23259516440783e-32 pua1 = -1.29304378590452e-37
+ ub1 = -7.02940198460963e-19 lub1 = -6.59229184468015e-24 wub1 = -4.13739827088341e-25 pub1 = 1.60737715953907e-30
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.84 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 4.2e-07 wmax = 7.0e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.014/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.785125784113331+0*(0.0/sqrt(l*w*mult))} lvth0 = -1.03594088297963e-08 wvth0 = -8.39141269016767e-08 pvth0 = 3.48291868541498e-14
+ k1 = 0.497655085274753 lk1 = 2.36596683902553e-08 wk1 = 4.48033604707344e-08 pk1 = -1.70464598398219e-14
+ k2 = 0.0702199064989271 lk2 = -1.75745938240541e-08 wk2 = -2.51139968580604e-08 pk2 = 1.20126095440641e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -236372.308804546 lvsat = 0.242822488033737 wvsat = 0.177849941252199 pvsat = -1.37296366304338e-7
+ ua = 1.87432032167266e-09 lua = 5.14935174198012e-16 wua = 1.12966282324632e-16 pua = -3.71349497292918e-22
+ ub = -2.31241292833985e-18 lub = 6.92424386955123e-25 wub = 1.46207693643934e-24 pub = -4.60216221071e-31
+ uc = 2.09155568097343e-11 luc = -1.88986165374996e-17 wuc = -1.70845677273193e-17 puc = 1.36161886346369e-23
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.00788064141241716 lu0 = 4.26633182715858e-09 wu0 = 7.1198522053438e-09 pu0 = -3.39306304282815e-15
+ a0 = 0.17470039286999 la0 = 6.47228713960621e-07 wa0 = 4.06814931982673e-07 pa0 = -4.66319227206631e-13
+ keta = -0.0969405415269949 lketa = 2.90395043760681e-08 wketa = 4.01381088885463e-08 pketa = -1.5433375019861e-14
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.994532904747236 lags = -7.38104119382722e-08 wags = -4.04993130980897e-07 pags = 5.31793684557581e-14
+ b0 = -2.12696788091484e-10 lb0 = 3.46430777552264e-13 wb0 = 2.32020453297225e-14 pb0 = -1.64520421309707e-19
+ b1 = -1.94270322577978e-08 lb1 = 1.80941076194482e-14 wb1 = 1.39412496176484e-14 pb1 = -1.28446979045342e-20
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {0.0791519077363501+0*(0.009/sqrt(l*w*mult))} lvoff = -8.77740086969307e-08 wvoff = -1.1159321313868e-07 pvoff = 6.32399444300169e-14
+ nfactor = {3.83380790040082+0*(0.02/sqrt(l*w*mult))} lnfactor = -1.67893354037198e-06 wnfactor = -1.33374424304734e-06 pnfactor = 1.13330197586943e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.78658214285714e-05 wcit = -5.66721421778571e-12
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -0.84407236185013 leta0 = 4.29046952243206e-07 weta0 = 6.666037393393e-07 peta0 = -3.37835055692756e-13
+ etab = 3.14176156740699 letab = -2.78925254808397e-06 wetab = -2.26082747927338e-06 petab = 2.0044002251536e-12
+ dsub = 0.415559229958778 ldsub = -2.18206934584332e-08 wdsub = -7.17629416810199e-08 pdsub = 1.57215041470927e-14
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -1.18665190253864 lpclm = 2.36187922497336e-06 wpclm = 1.69848212791526e-06 ppclm = -1.70170091528415e-12
+ pdiblc1 = 0.262060013107683 lpdiblc1 = 4.27306727205415e-07 wpdiblc1 = 2.05021357028618e-07 ppdiblc1 = -3.07868514657321e-13
+ pdiblc2 = 0.0030323531631973 lpdiblc2 = 3.0814541360053e-10 wpdiblc2 = -7.2170979100377e-10 ppdiblc2 = -2.22014456463392e-16
+ pdiblcb = -0.025
+ drout = 1.39514150731259 ldrout = -1.48444500835112e-06 wdrout = -6.98367063454042e-07 pdrout = 1.06952184628687e-12
+ pscbe1 = 277475322.861226 lpscbe1 = -42.3561016103147 wpscbe1 = 0.476404896306917 ppscbe1 = 3.05169782248093e-5
+ pscbe2 = 1.43535083640913e-08 lpscbe2 = -3.72812782191195e-16 wpscbe2 = 1.15608200751272e-16 ppscbe2 = 2.68606390189805e-22
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -2.44240149173481e-06 lalpha0 = -1.25041697927142e-11 walpha0 = 1.75978812977404e-12 palpha0 = 9.00907927727349e-18
+ alpha1 = 2.57316428571429e-10 walpha1 = -1.13344284355714e-16
+ beta0 = -40.8896330535695 lbeta0 = -1.29640266360255e-05 wbeta0 = 3.1621866160234e-05 pbeta0 = 9.34039969488349e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -1.33543054854293e-07 lagidl = 4.88132857618441e-14 wagidl = 9.629198474135e-14 pagidl = -3.5169289005408e-20
+ bgidl = 478897210.634649 lbgidl = -566.660050121217 wbgidl = 395.981115298684 pbgidl = 0.000408270632871635
+ cgidl = 3812.55416991509 lcgidl = -0.0025026231685146 wcgidl = -0.00111268302213858 pcgidl = 9.90677273198574e-10
+ egidl = -0.973186614151596 legidl = 1.8695212625478e-06 wegidl = 1.35657475567679e-06 pegidl = -1.34696389636802e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.814786468548714 lkt1 = 1.36467250516983e-07 wkt1 = 1.20167315578789e-07 pkt1 = -9.83227434559796e-14
+ kt2 = -0.019032
+ at = -431235.571003014 lat = 0.436036024700526 wat = 0.338832711646013 pat = -3.19927080629841e-7
+ ute = -1.74574759991245 lute = 2.61912146184517e-07 wute = 2.13226102470521e-07 pute = -1.88704034555899e-13
+ ua1 = 5.524e-10
+ ub1 = -3.77179350228825e-18 lub1 = -8.07518711232227e-25 wub1 = 1.30331235889654e-25 pub1 = 5.81805926180864e-31
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.81e-6
+ sbref = 2.81e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.85 pmos
* DC IV MOS Parameters
+ lmin = 8.0e-07 lmax = 1e-06 wmin = 4.2e-07 wmax = 7.0e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.02/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.651950411941627+0*(0.0/sqrt(l*w*mult))} lvth0 = -1.28218947324893e-07 wvth0 = -1.50863441530272e-07 pvth0 = 9.40789955538834e-14
+ k1 = 0.218824805399636 lk1 = 2.70423071928334e-07 wk1 = 2.45696673496838e-07 pk1 = -1.94836037401357e-13
+ k2 = 0.144784436230099 lk2 = -8.35638298134927e-08 wk2 = -8.77191720689297e-08 pk2 = 6.74178765798074e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -36335.5058283233 lvsat = 0.0657909175837953 wvsat = 0.0799914236634577 pvsat = -5.069206753089e-8
+ ua = 1.39646758651042e-09 lua = 9.37832455552916e-16 wua = 4.55342046553045e-16 pua = -6.74350336756245e-22
+ ub = -1.24691194233201e-19 lub = -1.24369840912059e-24 wub = 2.84342753700375e-25 pub = 5.82072641982072e-31
+ uc = -7.59244198328845e-13 luc = 2.83473980631308e-19 wuc = -1.46817704822385e-18 puc = -2.04239034409128e-25
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.00954978955959312 lu0 = 2.78914406264863e-09 wu0 = 6.60874413510624e-09 pu0 = -2.94073495620826e-15
+ a0 = 1.61674676078799 la0 = -6.28975111414974e-07 wa0 = -6.32159287453099e-07 pa0 = 4.53167762122929e-13
+ keta = -0.155890405467301 lketa = 8.1209839213919e-08 wketa = 8.88131603815137e-08 pketa = -5.85105522158797e-14
+ a1 = 0.0
+ a2 = 0.5
+ ags = 2.40808886271936 lags = -1.32480036696381e-06 wags = -1.4234404089164e-06 pags = 9.54500117192291e-13
+ b0 = 1.73121270979144e-06 lb0 = -1.18587205014359e-12 wb0 = -7.19933636015647e-13 pb0 = 4.93150941002538e-19
+ b1 = 4.50640603229222e-09 lb1 = -3.08686560009001e-15 wb1 = -2.53380849581732e-15 pb1 = 1.73564615059238e-21
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0142679717336129+0*(0.009/sqrt(l*w*mult))} lvoff = -5.09788246541073e-09 wvoff = -4.42854978588841e-08 pvoff = 3.67295294597392e-15
+ nfactor = {2.83653233349679+0*(0.02/sqrt(l*w*mult))} lnfactor = -7.96349650039747e-07 wnfactor = -7.28435165625091e-07 pnfactor = 5.97606468896126e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.78658214285714e-05 wcit = -5.66721421778571e-12
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.732132266903211 leta0 = -9.65886263180357e-07 weta0 = -5.01473578506019e-07 peta0 = 6.95907530213763e-13
+ etab = -0.00582533353225601 letab = -3.6538786872394e-09 wetab = 1.06965767512099e-09 petab = 2.63256843985436e-15
+ dsub = 1.4732717112157 ldsub = -9.57890950808406e-07 wdsub = -8.33829976451897e-07 pdsub = 6.90147019584145e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.60045012466508 lpclm = -1.04692133591801e-07 wpclm = -3.09585863256645e-07 ppclm = 7.54292165630229e-14
+ pdiblc1 = 0.64295564319814 lpdiblc1 = 9.0215999053511e-08 wpdiblc1 = -6.94086119127349e-08 ppdiblc1 = -6.49993642940678e-14
+ pdiblc2 = 0.0320402684226463 lpdiblc2 = -2.53637145514355e-08 wpdiblc2 = -2.16215066246231e-08 ppdiblc2 = 1.82742012423056e-14
+ pdiblcb = -0.025
+ drout = -2.24936633399572 ldrout = 1.74092620866752e-06 wdrout = 1.92744981309882e-06 pdrout = -1.25431296037803e-12
+ pscbe1 = 229250872.456703 lpscbe1 = 0.322295875436339 wpscbe1 = 35.2214462704603 ppscbe1 = -2.32209666109527e-7
+ pscbe2 = 1.15453162440313e-08 lpscbe2 = 2.11242320310137e-15 wpscbe2 = 2.13887130856489e-15 ppscbe2 = -1.5219713439097e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -7.33287570019603e-05 lalpha0 = 5.02299004020578e-11 walpha0 = 5.28324148659144e-11 palpha0 = -3.6189940021077e-17
+ alpha1 = 7.96121263517858e-10 lalpha1 = -4.76839584903415e-16 walpha1 = -5.01545624666927e-16 palpha1 = 3.43556245168722e-22
+ beta0 = -256.030662201346 lbeta0 = 0.000177434708454611 wbeta0 = 0.000186627965686799 pbeta0 = -1.27839223355629e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 3.32783081772591e-06 lagidl = -3.01448528460227e-12 wagidl = -2.39791108291315e-12 pagidl = 2.17218795485349e-18
+ bgidl = -1186048097.4518 lbgidl = 906.808222808749 wbgidl = 1595.55090054065 pbgidl = -0.000653342629218585
+ cgidl = 26568.2465770692 lcgidl = -0.0226412971703839 wcgidl = -0.0184258433901663 pcgidl = 1.63127376331012e-8
+ egidl = 7.80039784253015 legidl = -5.89505711369326e-06 wegidl = -4.96467001518002e-06 pegidl = 4.2473061196164e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.543760738097502 lkt1 = -1.03389165803688e-07 wkt1 = -7.63367521200092e-08 pkt1 = 7.55823739371183e-14
+ kt2 = -0.019032
+ at = 237723.752703572 lat = -0.155989631983183 wat = -0.100309124933385 pat = 6.87112490337443e-8
+ ute = -1.34705075 lute = -9.09325725037502e-8
+ ua1 = 5.524e-10
+ ub1 = -4.68424917857142e-18 wub1 = 7.8774277627221e-25
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.41e-6
+ sbref = 2.41e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.86 pmos
* DC IV MOS Parameters
+ lmin = 6e-07 lmax = 8.0e-07 wmin = 4.2e-07 wmax = 7.0e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.02/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.799668659786421+0*(0.0/sqrt(l*w*mult))} lvth0 = -2.70326861424486e-08 wvth0 = -2.65394716218313e-08 pvth0 = 8.91769778645136e-15
+ k1 = 0.579524378108619 lk1 = 2.33456681205441e-08 wk1 = -3.31390106816388e-08 pk1 = -3.83498791752209e-15
+ k2 = 0.0169974197124571 lk2 = 3.96963756600958e-09 wk2 = 1.01388034111012e-08 pk2 = 3.85652665863668e-16
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 112940.561680881 lvsat = -0.0364624422796719 wvsat = -0.0232505818545855 pvsat = 2.0028190038942e-8
+ ua = 7.97861401266154e-09 lua = -3.57090493562847e-15 wua = -2.40481911743914e-15 pua = 1.28484575977259e-21
+ ub = -1.21090809023122e-17 lub = 6.96554861896501e-24 wub = 5.08422020764973e-24 pub = -2.70581941458597e-30
+ uc = -1.21038847909782e-12 luc = 5.92505557236652e-19 wuc = -1.0590960122273e-18 puc = -4.84457498661578e-25
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0147414914528048 lu0 = -7.67145775691921e-10 wu0 = 3.16871817453502e-09 pu0 = -5.8433437334678e-16
+ a0 = -0.247288809432805 la0 = 6.47879934008423e-07 wa0 = 5.86856261021791e-07 pa0 = -3.81851793504628e-13
+ keta = 0.256007691078017 lketa = -2.00938297429141e-07 wketa = -1.37123763401597e-07 pketa = 9.62551108909323e-14
+ a1 = 0.0
+ a2 = 0.5
+ ags = -2.67839766625433 lags = 2.15941747295052e-06 wags = 1.33034215164695e-06 pags = -9.31827167880801e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {0.170334511274845+0*(0.009/sqrt(l*w*mult))} lvoff = -1.31549660313789e-07 wvoff = -1.22142619602204e-07 pvoff = 5.70046920545393e-14
+ nfactor = {3.17742468383073+0*(0.02/sqrt(l*w*mult))} lnfactor = -1.02985920555674e-06 wnfactor = 1.5348021934768e-07 pnfactor = -6.50116023329761e-15
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 6.81395370660714e-05 lcit = -3.44372438431093e-11 wcit = -3.31529198133355e-11 pcit = 1.88275709044236e-17
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -2.09186915780809 leta0 = 9.68540592739759e-07 weta0 = 1.55978567264891e-06 peta0 = -7.16044750531105e-13
+ etab = -0.175160371989742 letab = 1.12339775980946e-07 wetab = 1.15489282446556e-07 petab = -7.57443024304546e-14
+ dsub = -0.433924807584514 ldsub = 3.48529128587149e-07 wdsub = 5.84734669875514e-07 pdsub = -2.815626703269e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.5449559254212 lpclm = -6.66788845807383e-08 wpclm = -3.54479779116864e-07 ppclm = 1.06181324457692e-13
+ pdiblc1 = 0.263159881210096 lpdiblc1 = 3.50374197036511e-07 wpdiblc1 = 1.117878239989e-07 ppdiblc1 = -1.89118016911359e-13
+ pdiblc2 = -0.0330844521322543 lpdiblc2 = 1.92463934050686e-08 wpdiblc2 = 2.09061951744854e-08 ppdiblc2 = -1.08570618515748e-14
+ pdiblcb = -0.025
+ drout = -2.49485896086491 ldrout = 1.90908743060979e-06 wdrout = 1.10270152213474e-06 pdrout = -6.89364504809095e-13
+ pscbe1 = -240388597.390534 lpscbe1 = 322.022984523444 wpscbe1 = 160.67509849656 ppscbe1 = -8.61673341727269e-5
+ pscbe2 = 1.24158860867541e-08 lpscbe2 = 1.51608721368549e-15 wpscbe2 = 1.57125104241236e-15 ppscbe2 = -1.13315429969656e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -0.000138104160036267 lalpha0 = 9.4600727603543e-11 walpha0 = 3.96314739839897e-11 palpha0 = -2.7147361521663e-17
+ alpha1 = 3.424975e-10 lalpha1 = -1.661095750125e-16
+ beta0 = -126.585760989417 lbeta0 = 8.87655983489454e-05 wbeta0 = 1.21224027901131e-05 pbeta0 = -8.30378529921355e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -3.55107824172568e-06 lagidl = 1.69753302657677e-12 wagidl = 2.50825202158562e-12 pagidl = -1.18850924091265e-18
+ bgidl = -4358412478.22866 lbgidl = 3079.86196181899 wbgidl = 2636.86728873228 pbgidl = -0.00136663914854791
+ cgidl = -19923.2310121744 lcgidl = 0.00920513252085995 wcgidl = 0.0154096693061726 pcgidl = -6.86441938632743e-9
+ egidl = -3.59907497203189 legidl = 1.91352476691767e-06 wegidl = 3.17232994031427e-06 pegidl = -1.32649816489741e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.915888849983927 lkt1 = 1.51516730197955e-07 wkt1 = 1.16460402093364e-07 pkt1 = -5.6482712713271e-14
+ kt2 = -0.019032
+ at = 10000.0
+ ute = -1.434413128625 lute = -3.10897799575173e-08 wute = -2.74857055955498e-07 pute = 1.88275709044236e-13
+ ua1 = 5.5336999e-10 lua1 = -6.64438300049995e-19
+ ub1 = -1.15097030703777e-17 lub1 = 4.67540178861782e-24 wub1 = 2.69799931516293e-24 pub1 = -1.30851617785744e-30
+ uc1 = -5.5891912244259e-10 luc1 = 3.08055350277562e-16 wuc1 = 1.98094977368247e-16 puc1 = -1.35694069022362e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.02e-6
+ sbref = 2.01e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.87 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 6e-07 wmin = 4.2e-07 wmax = 7.0e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 5.75025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.0243e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.12565e-08+0*(1.12565e-08*(0.02/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.66132402464709+0*(0.0/sqrt(l*w*mult))} lvth0 = -9.41291424618487e-08 wvth0 = -1.69318882941004e-07 pvth0 = 7.81649983791931e-14
+ k1 = 0.826407699858027 lk1 = -9.63915085113091e-08 wk1 = -7.75870640392447e-08 pk1 = 1.772209572065e-14
+ k2 = -0.085811982941058 lk2 = 5.38316838059512e-08 wk2 = 2.13225845921401e-08 pk2 = -5.03842528803432e-15
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -41105.6111321819 lvsat = 0.0382491813037994 wvsat = 0.0440653426053009 pvsat = -1.26196967444805e-8
+ ua = -3.27613420905325e-10 lua = 4.5757383851429e-16 wua = -1.61731726111675e-15 pua = 9.02911296965506e-22
+ ub = 2.42541459137971e-18 lub = -8.36090229981201e-26 wub = 4.3766248872509e-24 pub = -2.36263922216914e-30
+ uc = 7.78934418710216e-12 luc = -3.77231978720701e-18 wuc = -1.43832557706784e-18 puc = -3.00533055861744e-25
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0134414070817505 lu0 = -1.36611356152461e-10 wu0 = 2.44031682675834e-09 pu0 = -2.3106336168182e-16
+ a0 = -1.33901481309204 la0 = 1.17736158715313e-06 wa0 = 1.90330420511671e-06 pa0 = -1.02032246415094e-12
+ keta = -0.346879758894143 lketa = 9.1459101370107e-08 wketa = 1.26887546395459e-07 pketa = -3.17890543040911e-14
+ a1 = 0.0
+ a2 = 0.5
+ ags = -1.04651800430356 lags = 1.36796399630271e-06 wags = 1.3440351556789e-06 pags = -9.38468206371279e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {0.000382925743880325+0*(0.009/sqrt(l*w*mult))} lvoff = -4.91239910891991e-08 wvoff = -9.98508229506505e-08 pvoff = 4.61932821375191e-14
+ nfactor = {-2.44732519317578+0*(0.02/sqrt(l*w*mult))} lnfactor = 1.69811636104203e-06 wnfactor = -3.90808849375137e-09 pnfactor = 6.98313821282579e-14
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -5.23985906375e-05 lcit = 2.40231454024843e-11 wcit = 2.74857055955498e-11 pcit = -1.05818592257587e-17
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -1.10978136355185 leta0 = 4.92232922964457e-07 weta0 = 6.83386611866359e-07 peta0 = -2.90995588046874e-13
+ etab = 0.187927043245021 letab = -6.37558049708374e-08 wetab = -1.23270764577949e-07 petab = 4.0053126576195e-14
+ dsub = 0.404641838205281 ldsub = -5.81715017876722e-08 wdsub = -2.44206984306676e-08 pdsub = 1.38746375247563e-14
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 3.14630210830381 lpclm = -8.43323776547887e-07 wpclm = -8.88671968755207e-07 ppclm = 3.65261865471341e-13
+ pdiblc1 = 5.34562888937674 lpdiblc1 = -2.11459785957927e-06 wpdiblc1 = -2.25702898951189e-06 ppdiblc1 = 9.59746293557309e-13
+ pdiblc2 = 0.0375648513101968 lpdiblc2 = -1.5018165518003e-08 wpdiblc2 = -2.14592888164833e-08 ppdiblc2 = 9.68998605662507e-15
+ pdiblcb = -0.025
+ drout = 2.09056696400399 ldrout = -3.14821215822001e-07 wdrout = -7.8878768868693e-07 pdrout = 2.27998304993363e-13
+ pscbe1 = 286050046.447241 lpscbe1 = 66.7028744553425 wpscbe1 = 82.0993462354131 ppscbe1 = -4.80584872048319e-5
+ pscbe2 = 1.8374315413026e-08 lpscbe2 = -1.37372121740978e-15 wpscbe2 = -3.53143981909769e-15 ppscbe2 = 1.34162525468151e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.000150161416231063 lalpha0 = -4.52066355582308e-11 walpha0 = -4.23609233131291e-11 palpha0 = 1.26185412054531e-17
+ alpha1 = 0.0
+ beta0 = 74.893242785407 lbeta0 = -8.95071108682511e-06 wbeta0 = -1.03120799034637e-05 pbeta0 = 2.57682663475772e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -3.25133577033436e-07 lagidl = 1.32965993924356e-13 wagidl = 2.43847609172142e-13 pagidl = -9.02844229141734e-20
+ bgidl = 2105848674.51472 lbgidl = -55.2723759557775 wbgidl = -383.746333699357 pbgidl = 9.83433552633264e-5
+ cgidl = -8245.68534569617 lcgidl = 0.00354158126034636 wcgidl = 0.00640633624895125 pcgidl = -2.49784787024035e-9
+ egidl = -0.54482369079307 legidl = 4.32228166773245e-07 wegidl = 1.14590243524599e-06 pegidl = -3.43690957076816e-13
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.436288853841787 lkt1 = -8.10868699310028e-08 wkt1 = 4.36369827555309e-09 pkt1 = -2.11637184515185e-15
+ kt2 = -0.019032
+ at = 107985.599943214 lat = -0.0475225260444592 wat = -0.0567280775821867 pat = 2.75128339869727e-8
+ ute = -1.95123068508915 lute = 2.19564150839808e-07 wute = 5.18295484327017e-07 pute = -1.96399307230081e-13
+ ua1 = 5.52e-10
+ ub1 = -6.15642282890016e-20 lub1 = -8.76888309100974e-25 wub1 = 9.40813348209191e-25 pub1 = -4.56289769814716e-31
+ uc1 = 1.20029455138944e-09 luc1 = -5.45154485462604e-16 wuc1 = -6.91629782784522e-16 puc1 = 2.9581799102793e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.52493723e-10
+ cgso = 1.52493723e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.7168565e-12
+ cgdl = 7.7168565e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 5.71105e-8
+ dwc = -2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007398371535
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.513752158e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.4070604e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 1.81e-6
+ sbref = 1.81e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.ends sky130_fd_pr__pfet_g5v0d10v5
