* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
.subckt  sky130_fd_pr__pfet_g5v0d10v5 d g s b
+ 
.param  l = 1 w = 1 ad = 0 as = 0 pd = 0 ps = 0 nrd = 0 nrs = 0 sa = 0 sb = 0 sd = 0 mult = 1 nf = 1.0
msky130_fd_pr__pfet_g5v0d10v5 d g s b sky130_fd_pr__pfet_g5v0d10v5__model l = {l} w = {w} ad = {ad} as = {as} pd = {pd} ps = {ps} nrd = {nrd} nrs = {nrs} sa = {sa} sb = {sb} sd = {sd} nf = {nf}
.model sky130_fd_pr__pfet_g5v0d10v5__model.0 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 2.0e-05 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.964555+0*(0.0/sqrt(l*w*mult))}
+ k1 = 0.59521
+ k2 = 0.02039548
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200000.0
+ ua = 2.7054732e-9
+ ub = -5.157e-20
+ uc = -3.9972e-11
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0209529
+ a0 = 0.8941253
+ keta = -0.0079259
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.1386898
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.093204657+0*(0.009/sqrt(l*w*mult))}
+ nfactor = {1.79934+0*(0.02/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.080000000000001
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.08353125
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0029407877
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 333712830.0
+ pscbe2 = 1.5000958e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 5.0667189e-5
+ alpha1 = 0.0
+ beta0 = 38.266046
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 7.3657e-9
+ bgidl = 1704700000.0
+ cgidl = 700.0
+ egidl = 0.69350825
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.57573
+ kt2 = -0.019032
+ at = 430000.0
+ ute = -1.3864
+ ua1 = 7.0656e-10
+ ub1 = -3.145e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.1 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 2.0e-05 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.964555+0*(0.0/sqrt(l*w*mult))}
+ k1 = 0.59521
+ k2 = 0.02039548
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200000.0
+ ua = 2.7054732e-9
+ ub = -5.157e-20
+ uc = -3.9972e-11
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0209529
+ a0 = 0.8941253
+ keta = -0.0079259
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.1386898
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.093204657+0*(0.009/sqrt(l*w*mult))}
+ nfactor = {1.79934+0*(0.02/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.080000000000001
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.08353125
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0029407877
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 333712830.0
+ pscbe2 = 1.5000958e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 5.0667189e-5
+ alpha1 = 0.0
+ beta0 = 38.266046
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 7.3657e-9
+ bgidl = 1704700000.0
+ cgidl = 700.0
+ egidl = 0.69350825
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.57573
+ kt2 = -0.019032
+ at = 430000.0
+ ute = -1.3864
+ ua1 = 7.0656e-10
+ ub1 = -3.145e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.2 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 2.0e-05 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.9708996575+0*(0.0/sqrt(l*w*mult))} lvth0 = 4.99616399495017e-8
+ k1 = 0.6040731475 lk1 = -6.97937413035002e-8
+ k2 = 0.017946422832 lk2 = 1.92853455751328e-8
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 296855.3135 lvsat = -0.7626968516871
+ ua = 2.452507249685e-09 lua = 1.9920056723505e-15
+ ub = 2.05160996e-19 lub = -2.0216539011016e-24 wub = -3.67341984631965e-40 pub = 4.20389539297445e-45
+ uc = -5.147278145e-11 luc = 9.05640536061701e-17
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.020337710385 lu0 = 4.844372142279e-9
+ a0 = 0.913768069025 la0 = -1.54678948964264e-7
+ keta = -0.004983044435 lketa = -2.3173810432149e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.113393989575 lags = 1.99194388772705e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0947625464815+0*(0.009/sqrt(l*w*mult))} lvoff = 1.22677565110199e-8
+ nfactor = {1.8039023415+0*(0.02/sqrt(l*w*mult))} lnfactor = -3.5926614375899e-8
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.080000000000001
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.641832441643 lpclm = 5.71194892621197e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 0.004539823205605 lpdiblc2 = -1.25917649924371e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 560098762.7795 lpscbe1 = -1782.69866626545
+ pscbe2 = -1.50486592213e-08 lpscbe2 = 2.36628715770849e-13
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 7.7909598465e-05 lalpha0 = -2.14523077573089e-10
+ alpha1 = 0.0
+ beta0 = 39.13253926505 lbeta0 = -6.82328786496275e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 6.546125235e-09 lagidl = 6.453823444469e-15
+ bgidl = 1480360660 lbgidl = 1766.582566764
+ cgidl = 930.5387 lcgidl = -0.00181540004702
+ egidl = 1.2047468705955 legidl = -4.02579964174133e-6
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.5851549645 lkt1 = 7.42178254517005e-8
+ kt2 = -0.019032
+ at = 670893.5685 lat = -1.8969404945101
+ ute = -1.222020095 lute = -1.294425999913e-6
+ ua1 = 1.3695660536e-09 lua1 = -5.22090746967856e-15
+ ub1 = -2.61514845e-18 lub1 = -4.17236901563001e-24
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.3 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 2.0e-05 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.9431553561+0*(0.0/sqrt(l*w*mult))} lvth0 = -5.75364302549401e-8
+ k1 = 0.602294036 lk1 = -6.29003958856002e-8
+ k2 = 0.023211373013 lk2 = -1.1142303961698e-9
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 84825.74 lvsat = 0.058832933796
+ ua = 3.31328698619e-09 lua = -1.34317149471177e-15
+ ub = -1.239166271e-18 lub = 3.5745365276166e-24
+ uc = -5.44361927e-11 luc = 1.0204608683542e-16
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.02075923934 lu0 = 3.21111605323601e-9
+ a0 = 0.825992817278 la0 = 1.85415041454661e-7
+ keta = -0.0051939812 lketa = -2.235651484248e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.13791869307 lags = 1.04170972610978e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0645862731911+0*(0.009/sqrt(l*w*mult))} lvoff = -1.04653231979964e-7
+ nfactor = {2.231805466+0*(0.02/sqrt(l*w*mult))} lnfactor = -1.6938800605636e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.020200260000001 leta0 = 2.31700072604e-7
+ etab = -0.1214502716 letab = 1.9934922234136e-7
+ dsub = 0.810118505 ldsub = -9.69109159473e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.044838468325 lpclm = -8.23226181550045e-7
+ pdiblc1 = 0.57808555402 lpdiblc1 = -7.28756287605892e-7
+ pdiblc2 = -0.0010893622944 lpdiblc2 = 9.21907714588224e-9
+ pdiblcb = 0.16246 lpdiblcb = -7.26332516e-07 wpdiblcb = 2.11758236813575e-22
+ drout = 0.147588 ldrout = 1.5979315352e-6
+ pscbe1 = -151521249.434 lpscbe1 = 974.544233056976 ppscbe1 = 1.73472347597681e-18
+ pscbe2 = 7.55293005675e-08 lpscbe2 = -1.14324647226835e-13
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 4.36726325897e-05 lalpha0 = -8.18685295926516e-11
+ alpha1 = -9.373e-11 lalpha1 = 3.63166258e-16
+ beta0 = 69.5879243857 lbeta0 = -0.000124825723053433 pbeta0 = 4.13590306276514e-25
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 9.17928106e-09 lagidl = -3.748602115076e-15
+ bgidl = 2607594260 lbgidl = -2600.996739796
+ cgidl = 455.860685 lcgidl = 2.37873898990002e-5
+ egidl = -1.553543708466 legidl = 6.66147303589036e-06 wegidl = -3.3881317890172e-21 pegidl = -6.46234853557053e-27
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.5669373 lkt1 = 3.6316625799996e-9
+ kt2 = -0.019032
+ at = 209907.023 lat = -0.1108020253158
+ ute = -1.70241253 lute = 5.66902528738e-7
+ ua1 = -4.749579392e-10 lua1 = 1.92588519282432e-15 wua1 = 7.88860905221012e-31 pua1 = -2.63310734584192e-36
+ ub1 = -3.71946289e-18 lub1 = 1.06407713594004e-25
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.4 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 2.0e-05 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.9966077158+0*(0.0/sqrt(l*w*mult))} lvth0 = 4.26653632386798e-8
+ k1 = 0.55942551 lk1 = 1.74609429539997e-8
+ k2 = 0.017219824654 lk2 = 1.01175261576116e-8
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 175963.5466 lvsat = -0.11201399845636
+ ua = 3.424749578434e-09 lua = -1.55211927013238e-15
+ ub = 6.4325866e-19 lub = 4.57427519639998e-26
+ uc = 5.12043316e-13 luc = -9.598764001736e-19
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.02566702634 lu0 = -5.989021456964e-9
+ a0 = 1.000482195724 la0 = -1.4168274738021e-7
+ keta = 0.0419609792 lketa = -1.1075320360832e-07 pketa = 2.01948391736579e-28
+ a1 = 0.0
+ a2 = 0.5
+ ags = -0.29536367256 lags = 9.16402095220976e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1577214518922+0*(0.009/sqrt(l*w*mult))} lvoff = 6.99379740131181e-8
+ nfactor = {1.088455902+0*(0.02/sqrt(l*w*mult))} lnfactor = 4.49443032110801e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.4373e-05 lcit = -8.1976258e-12
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.269542430581401 leta0 = -2.35716760367893e-7
+ etab = -0.0283214568 letab = 2.476994611728e-8
+ dsub = 0.0736166540000002 ldsub = 4.115372104116e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.083196751172 lpclm = 9.79467381424969e-7
+ pdiblc1 = 0.00549710252000002 lpdiblc1 = 3.44618023576008e-7
+ pdiblc2 = 0.00585964945018 lpdiblc2 = -3.80754027050743e-9
+ pdiblcb = -0.39992 lpdiblcb = 3.27905032e-7
+ drout = 1.515411042014 ldrout = -9.66189539359445e-07 wdrout = 6.7762635780344e-21
+ pscbe1 = 428577028.488 lpscbe1 = -112.907998735605
+ pscbe2 = 1.45331535696e-08 lpscbe2 = 1.87299354278389e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -5.93092031506e-05 lalpha0 = 1.11181219686115e-10 walpha0 = 6.58698855859545e-27 palpha0 = -1.82584177258986e-31
+ alpha1 = 1.8746e-10 lalpha1 = -1.63952516e-16
+ beta0 = -38.239948205 lbeta0 = 7.7308406905093e-05 pbeta0 = 5.16987882845642e-26
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 3.96946816e-09 lagidl = 6.017713147264e-15
+ bgidl = 869210480 lbgidl = 657.777494192
+ cgidl = 440.624022 lcgidl = 5.23500383587999e-5
+ egidl = 3.067904826664 legidl = -2.00189438806434e-6
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.50272848 lkt1 = -1.16734191392e-7
+ kt2 = -0.019032
+ at = 256626.6 lat = -0.19838254436
+ ute = -1.21904526 lute = -3.39217755604e-7
+ ua1 = 6.68354468e-10 lua1 = -2.173682457128e-16
+ ub1 = -3.53701998e-18 lub1 = -2.35599765492001e-25
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.81e-6
+ sbref = 2.81e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.5 pmos
* DC IV MOS Parameters
+ lmin = 8.0e-07 lmax = 1e-06 wmin = 2.0e-05 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.053103076+0*(0.0/sqrt(l*w*mult))} lvth0 = 9.20762052695999e-8
+ k1 = 0.589711379999999 lk1 = -9.02707894799971e-9
+ k2 = 0.0122474826 lk2 = 1.446633651804e-8
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 12212.779 lvsat = 0.0312024228866
+ ua = -7.00597444169999e-10 lua = 2.05590923583708e-15
+ ub = 3.95360816e-18 lub = -2.849488920736e-24 wub = 1.17549435082229e-38
+ uc = 5.75692682e-12 luc = -5.547051512772e-18 puc = 5.87747175411144e-39
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0203449079 lu0 = -1.33429666934e-9
+ a0 = 0.821535675 la0 = 1.48238796449997e-8
+ keta = -0.150384786 lketa = 5.74724026356e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.858047376 lags = -9.23712078496003e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0943996895959999+0*(0.009/sqrt(l*w*mult))} lvoff = 1.45567607088615e-8
+ nfactor = {0.732679410000001+0*(0.02/sqrt(l*w*mult))} lnfactor = 7.60605152014001e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -1.1865e-05 lcit = 1.4750129e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -6.676430499899e-05 leta0 = 8.3441479753e-11
+ etab = 0.00071767321 letab = -6.27676989466e-10
+ dsub = 1.45264382 ldsub = -7.94559948971999e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.98189989655 lpclm = -6.8113838952263e-7
+ pdiblc1 = 0.20581194057 lpdiblc1 = 1.69422666217478e-7
+ pdiblc2 = -0.0319025077049 lpdiblc2 = 2.92192423773255e-08 ppdiblc2 = -5.04870979341448e-29
+ pdiblcb = -0.025
+ drout = 0.33949907438 ldrout = 6.22630675332523e-8
+ pscbe1 = -39572648.0999999 lpscbe1 = 296.53570840826
+ pscbe2 = 1.8099436842e-08 lpscbe2 = -3.1003414146132e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.00023839585627 lalpha0 = -1.49191625283142e-10
+ alpha1 = 0.0
+ beta0 = 66.364220735 lbeta0 = -1.4178399249831e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 9.12977e-09 lagidl = 1.50451315800001e-15
+ bgidl = 993921999.999999 lbgidl = 548.7047988
+ cgidl = 434.63904 lcgidl = 5.75845036159999e-5
+ egidl = 1.78393816687 legidl = -8.78937147408502e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.6115771 lkt1 = -2.15351883400002e-8
+ kt2 = -0.019032
+ at = 45990.4 lat = -0.01416012384
+ ute = -2.0356083 lute = 3.7494827918e-7
+ ua1 = -2.73723399999993e-11 lua1 = 3.91114420564e-16
+ ub1 = -4.5332815e-18 lub1 = 6.35730559899999e-25
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.41e-6
+ sbref = 2.41e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.6 pmos
* DC IV MOS Parameters
+ lmin = 6e-07 lmax = 8.0e-07 wmin = 2.0e-05 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.866730167+0*(0.0/sqrt(l*w*mult))} lvth0 = -3.36509591417997e-8
+ k1 = 0.59315457 lk1 = -1.1349854922e-8
+ k2 = 0.0156090654 lk2 = 1.219861276116e-8
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 59706.6044 lvsat = -0.000836911728240006
+ ua = -1.7341739129e-09 lua = 2.75315992164234e-15
+ ub = 2.4292250742e-18 lub = -1.82114009105532e-24 pub = 2.80259692864963e-45
+ uc = 2.4254276e-12 luc = -3.29962213896e-18
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0075359161 lu0 = 7.30664919894001e-9
+ a0 = 0.93256869 la0 = -6.0078992274e-8
+ keta = 0.010069695 lketa = -5.0770190247e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = -0.53391224 lags = 8.46644749104e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {0.00559779755700002+0*(0.009/sqrt(l*w*mult))} lvoff = -5.29015441245522e-8
+ nfactor = {1.7678603+0*(0.02/sqrt(l*w*mult))} lnfactor = 6.22721236199998e-8
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -0.056074191601999 leta0 = 3.78660519343092e-08 weta0 = 2.23338765389317e-23 peta0 = -5.28536806498078e-29
+ etab = -0.00071767321 letab = 3.40607705466e-10
+ dsub = 0.19513736522 ldsub = 5.3753905422588e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.27276388295 lpclm = 4.7184476525193e-7
+ pdiblc1 = 0.19544523505 lpdiblc1 = 1.7641604576127e-7
+ pdiblc2 = 0.0256746597612 lpdiblc2 = -9.62231479530552e-9
+ pdiblcb = -0.025
+ drout = -0.65870811482 ldrout = 7.35653637367572e-7
+ pscbe1 = 430031833.72 lpscbe1 = -20.2594750275119
+ pscbe2 = 1.0746893781e-08 lpscbe2 = 1.8596841343374e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -0.000112188837415 lalpha0 = 8.7312809076759e-11 walpha0 = 2.06795153138257e-25 palpha0 = 9.86076131526265e-32
+ alpha1 = 0.0
+ beta0 = 27.750617018 lbeta0 = 1.18703378176572e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 2.28427097e-08 lagidl = -7.74623596362e-15
+ bgidl = 2044837300.0 lbgidl = -160.24266258
+ cgidl = 1208.17 lcgidl = -0.000464239482
+ egidl = -0.1972262296 legidl = 4.5755635445016e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.70287246 lkt1 = 4.00526615159997e-8
+ kt2 = -0.019032
+ at = 41611 lat = -0.0112057806
+ ute = -1.6043825 lute = 8.40433545e-8
+ ua1 = 5.533492e-10 lua1 = -6.40330320000131e-19
+ ub1 = -4.2831041e-18 lub1 = 4.6696088586e-25
+ uc1 = -2.69861592e-10 luc1 = 1.083823099632e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.02e-6
+ sbref = 2.01e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.7 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 6e-07 wmin = 2.0e-05 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.02/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.845928173999999+0*(0.0/sqrt(l*w*mult))} lvth0 = -4.35235850196003e-8
+ k1 = 0.4613552 lk1 = 5.12021260800003e-8
+ k2 = 0.037165178 lk2 = 1.96808172119999e-9
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 38567.015 lvsat = 0.00919593740100003
+ ua = 1.121182010942e-08 lua = -3.39100884135074e-15
+ ub = -7.30555818840001e-18 lub = 2.79898804537464e-24
+ uc = -1.700643e-12 luc = -1.3413890322e-18
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.036021697 lu0 = -6.2127024162e-9
+ a0 = 0.23036964 la0 = 2.73184676856001e-7
+ keta = -0.13824211 lketa = 1.9618592406e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 1.25
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.12209155362+0*(0.009/sqrt(l*w*mult))} lvoff = 7.699821944052e-9
+ nfactor = {1.32304758+0*(0.02/sqrt(l*w*mult))} lnfactor = 2.73380240532001e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 2.873e-05 lcit = -8.88925800000001e-12
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -0.187353623999999 leta0 = 1.001712705504e-7
+ etab = 0.0144232238 letab = -6.84526201548001e-9
+ dsub = 0.41601716956 ldsub = -5.10756497171761e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.006081441 lpclm = 1.238122522014e-7
+ pdiblc1 = 1.59030588952 lpdiblc1 = -4.85584820850193e-7
+ pdiblc2 = 0.00764468105400001 lpdiblc2 = -1.0652869008684e-9
+ pdiblcb = -0.025
+ drout = 0.86038901644 ldrout = 1.46901388715762e-8
+ pscbe1 = 479887042.4 lpscbe1 = -43.9207570670401
+ pscbe2 = 1.5334308648e-08 lpscbe2 = -3.17502961540804e-16
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -2.31891527040001e-05 lalpha0 = 4.50735587129184e-11
+ alpha1 = 0.0
+ beta0 = 45.559628338 lbeta0 = 3.4181810451852e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -2.10753074e-08 lagidl = 1.309725495204e-14
+ bgidl = 2054454200.0 lbgidl = -164.80684332
+ cgidl = -2189.916 lcgidl = 0.0011484921336 wcgidl = -3.46944695195361e-18 pcgidl = -1.65436122510606e-24
+ egidl = 1.1474310464 legidl = -1.8061798873944e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.63721 lkt1 = 8.88925800000003e-9
+ kt2 = -0.019032
+ at = 18000.0
+ ute = -1.6329554 lute = 9.760405284e-8
+ ua1 = 5.52e-10
+ ub1 = -7.56664320000001e-18 lub1 = 2.02532854272e-24
+ uc1 = -4.1496e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 1.81e-6
+ sbref = 1.81e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.8 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 1.5e-05 wmax = 2.0e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.964555+0*(0.0/sqrt(l*w*mult))}
+ k1 = 0.59521
+ k2 = 0.02039548
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200000.0
+ ua = 2.7054732e-9
+ ub = -5.157e-20
+ uc = -3.9972e-11
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0209529
+ a0 = 0.8941253
+ keta = -0.0079259
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.1386898
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.093204657+0*(0.009/sqrt(l*w*mult))}
+ nfactor = {1.79934+0*(0.02/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.080000000000001
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.08353125
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0029407877
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 333712830.0
+ pscbe2 = 1.5000958e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 5.0667189e-5
+ alpha1 = 0.0
+ beta0 = 38.266046
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 7.3657e-9
+ bgidl = 1704700000.0
+ cgidl = 700.0
+ egidl = 0.69350825
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.57573
+ kt2 = -0.019032
+ at = 430000.0
+ ute = -1.3864
+ ua1 = 7.0656e-10
+ ub1 = -3.145e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.9 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 1.5e-05 wmax = 2.0e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.964555+0*(0.0/sqrt(l*w*mult))}
+ k1 = 0.59521
+ k2 = 0.02039548
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200000.0
+ ua = 2.7054732e-9
+ ub = -5.157e-20
+ uc = -3.9972e-11
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0209529
+ a0 = 0.8941253
+ keta = -0.0079259
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.1386898
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.093204657+0*(0.009/sqrt(l*w*mult))}
+ nfactor = {1.79934+0*(0.02/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.080000000000001
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.08353125
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0029407877
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 333712830.0
+ pscbe2 = 1.5000958e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 5.0667189e-5
+ alpha1 = 0.0
+ beta0 = 38.266046
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 7.3657e-9
+ bgidl = 1704700000.0
+ cgidl = 700.0
+ egidl = 0.69350825
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.57573
+ kt2 = -0.019032
+ at = 430000.0
+ ute = -1.3864
+ ua1 = 7.0656e-10
+ ub1 = -3.145e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.10 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 1.5e-05 wmax = 2.0e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.9708996575+0*(0.0/sqrt(l*w*mult))} lvth0 = 4.99616399495e-8
+ k1 = 0.604073147499999 lk1 = -6.9793741303501e-8
+ k2 = 0.017946422832 lk2 = 1.92853455751329e-8
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 296855.3135 lvsat = -0.7626968516871
+ ua = 2.452507249685e-09 lua = 1.99200567235049e-15
+ ub = 2.05160996e-19 lub = -2.0216539011016e-24 pub = -8.4077907859489e-45
+ uc = -5.14727814500001e-11 luc = 9.056405360617e-17
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.020337710385 lu0 = 4.84437214227905e-9
+ a0 = 0.913768069025001 la0 = -1.54678948964262e-7
+ keta = -0.00498304443499999 lketa = -2.3173810432149e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.113393989575 lags = 1.99194388772706e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0947625464815+0*(0.009/sqrt(l*w*mult))} lvoff = 1.22677565110199e-8
+ nfactor = {1.8039023415+0*(0.02/sqrt(l*w*mult))} lnfactor = -3.59266143758956e-8
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.080000000000001
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.641832441643 lpclm = 5.71194892621197e-06 wpclm = 1.6940658945086e-21 ppclm = -6.46234853557053e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 0.004539823205605 lpdiblc2 = -1.25917649924371e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 560098762.7795 lpscbe1 = -1782.69866626545
+ pscbe2 = -1.50486592213e-08 lpscbe2 = 2.36628715770849e-13 ppscbe2 = 7.70371977754894e-34
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 7.7909598465e-05 lalpha0 = -2.14523077573089e-10
+ alpha1 = 0.0
+ beta0 = 39.13253926505 lbeta0 = -6.82328786496275e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 6.546125235e-09 lagidl = 6.45382344446899e-15
+ bgidl = 1480360660.0 lbgidl = 1766.582566764
+ cgidl = 930.5387 lcgidl = -0.00181540004702
+ egidl = 1.2047468705955 legidl = -4.02579964174132e-06 pegidl = -5.16987882845642e-26
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.5851549645 lkt1 = 7.42178254516996e-8
+ kt2 = -0.019032
+ at = 670893.5685 lat = -1.8969404945101
+ ute = -1.222020095 lute = -1.294425999913e-6
+ ua1 = 1.3695660536e-09 lua1 = -5.22090746967856e-15
+ ub1 = -2.61514845e-18 lub1 = -4.17236901563e-24
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.11 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 1.5e-05 wmax = 2.0e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.9431553561+0*(0.0/sqrt(l*w*mult))} lvth0 = -5.75364302549401e-8
+ k1 = 0.602294036 lk1 = -6.29003958856006e-8
+ k2 = 0.023211373013 lk2 = -1.11423039616984e-9
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 84825.7400000001 lvsat = 0.0588329337960001
+ ua = 3.31328698619e-09 lua = -1.34317149471177e-15
+ ub = -1.239166271e-18 lub = 3.5745365276166e-24 pub = 1.12103877145985e-44
+ uc = -5.44361927e-11 luc = 1.0204608683542e-16
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.02075923934 lu0 = 3.21111605323603e-9
+ a0 = 0.825992817278 la0 = 1.85415041454661e-7
+ keta = -0.0051939812 lketa = -2.235651484248e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.13791869307 lags = 1.04170972610978e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0645862731910999+0*(0.009/sqrt(l*w*mult))} lvoff = -1.04653231979964e-7
+ nfactor = {2.231805466+0*(0.02/sqrt(l*w*mult))} lnfactor = -1.6938800605636e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.0202002600000011 leta0 = 2.31700072604e-7
+ etab = -0.1214502716 letab = 1.9934922234136e-7
+ dsub = 0.810118505 ldsub = -9.69109159473001e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.044838468325 lpclm = -8.23226181550045e-7
+ pdiblc1 = 0.578085554019999 lpdiblc1 = -7.28756287605892e-7
+ pdiblc2 = -0.0010893622944 lpdiblc2 = 9.21907714588224e-09 ppdiblc2 = 5.04870979341448e-29
+ pdiblcb = 0.16246 lpdiblcb = -7.26332516e-07 wpdiblcb = 8.470329472543e-22 ppdiblcb = -1.61558713389263e-27
+ drout = 0.147588 ldrout = 1.5979315352e-6
+ pscbe1 = -151521249.434 lpscbe1 = 974.544233056976
+ pscbe2 = 7.55293005675e-08 lpscbe2 = -1.14324647226836e-13
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 4.36726325897e-05 lalpha0 = -8.18685295926517e-11
+ alpha1 = -9.37299999999999e-11 lalpha1 = 3.63166258e-16
+ beta0 = 69.5879243857 lbeta0 = -0.000124825723053433
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 9.17928105999999e-09 lagidl = -3.748602115076e-15
+ bgidl = 2607594260.0 lbgidl = -2600.996739796
+ cgidl = 455.860685 lcgidl = 2.37873898989993e-5
+ egidl = -1.553543708466 legidl = 6.66147303589036e-06 wegidl = 3.3881317890172e-21
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.566937299999999 lkt1 = 3.63166257999917e-9
+ kt2 = -0.019032
+ at = 209907.023 lat = -0.1108020253158
+ ute = -1.70241253 lute = 5.66902528738001e-7
+ ua1 = -4.749579392e-10 lua1 = 1.92588519282432e-15 wua1 = 1.18329135783152e-30 pua1 = 4.51389830715758e-36
+ ub1 = -3.71946289e-18 lub1 = 1.06407713594001e-25
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.12 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 1.5e-05 wmax = 2.0e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.996791869078143+0*(0.0/sqrt(l*w*mult))} lvth0 = 4.3010576973886e-08 wvth0 = 3.69039412670782e-09 pvth0 = -6.91801282992006e-15
+ k1 = 0.55942551 lk1 = 1.74609429539999e-8
+ k2 = 0.0159625839165107 lk2 = 1.24743496441091e-08 wk2 = 2.51948479021759e-08 pk2 = -4.72302618774187e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 175963.5466 lvsat = -0.11201399845636 wvsat = -1.77635683940025e-15
+ ua = 3.42652873586936e-09 lua = -1.55545447866069e-15 wua = -3.56539520564474e-17 pua = 6.68368985249868e-23
+ ub = 1.43532821690163e-18 lub = -1.43907083940379e-24 wub = -1.5872912338119e-23 pub = 2.97553614690378e-29
+ uc = 5.12043316e-13 luc = -9.59876400173601e-19
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0273694970888153 lu0 = -9.1804731226932e-09 wu0 = -3.41171665022266e-08 pu0 = 6.39560403250736e-14
+ a0 = 0.987370482320261 la0 = -1.17103529433562e-07 wa0 = 2.62756061821391e-07 pa0 = -4.92562513490391e-13
+ keta = 0.0419609792 lketa = -1.1075320360832e-7
+ a1 = 0.0
+ a2 = 0.5
+ ags = -0.316215085167952 lags = 9.55490153295843e-07 wags = 4.17858054975189e-07 pags = -7.83316709856488e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1577214518922+0*(0.009/sqrt(l*w*mult))} lvoff = 6.99379740131183e-8
+ nfactor = {1.25932383650498+0*(0.02/sqrt(l*w*mult))} lnfactor = 1.29134002087758e-07 wnfactor = -3.42415855042125e-06 pnfactor = 6.41892761861963e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.4373e-05 lcit = -8.1976258e-12
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.269577887979727 leta0 = -2.35783228806794e-07 weta0 = -7.10559029140184e-10 peta0 = 1.33201395602317e-15
+ etab = -0.0283214568 letab = 2.476994611728e-8
+ dsub = 0.0736166540000003 ldsub = 4.11537210411601e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.0831967511720002 lpclm = 9.7946738142497e-7
+ pdiblc1 = 0.00549710251999991 lpdiblc1 = 3.44618023576008e-7
+ pdiblc2 = 0.00585964945018 lpdiblc2 = -3.80754027050743e-9
+ pdiblcb = -0.39992 lpdiblcb = 3.27905032e-07 ppdiblcb = -3.23117426778526e-27
+ drout = 1.515411042014 ldrout = -9.66189539359445e-7
+ pscbe1 = 428577028.488 lpscbe1 = -112.907998735604
+ pscbe2 = 1.45331535696e-08 lpscbe2 = 1.87299354278452e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -5.93092031506e-05 lalpha0 = 1.11181219686115e-10 walpha0 = -1.49004780943576e-25 palpha0 = 1.53359694985679e-31
+ alpha1 = 1.8746e-10 lalpha1 = -1.63952516e-16
+ beta0 = -38.239948205 lbeta0 = 7.7308406905093e-05 wbeta0 = -1.0842021724855e-19 pbeta0 = -3.6189151799195e-25
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -2.61690537081875e-09 lagidl = 1.83645289681368e-14 wagidl = 1.31989581937407e-13 pagidl = -2.47427670299864e-19
+ bgidl = 1047049931.46323 lbgidl = 324.399658479026 wbgidl = -3563.86632807506 pbgidl = 0.00668082381860952
+ cgidl = 92.1007893099268 lcgidl = 0.000705691690359612 wcgidl = 0.0069843344843696 pcgidl = -1.30928334243993e-8
+ egidl = 3.067904826664 legidl = -2.00189438806434e-06 pegidl = -2.58493941422821e-26
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.5158822855816 lkt1 = -9.20760674487327e-08 wkt1 = 2.63599580478929e-07 pkt1 = -4.94143773565787e-13
+ kt2 = -0.019032
+ at = 261888.12223264 lat = -0.208245793937307 wat = -0.105439832191571 pat = 1.97657509426317e-7
+ ute = -1.21904526 lute = -3.39217755604001e-7
+ ua1 = 6.68354468e-10 lua1 = -2.173682457128e-16
+ ub1 = -3.53701998e-18 lub1 = -2.35599765492001e-25
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.81e-6
+ sbref = 2.81e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.13 pmos
* DC IV MOS Parameters
+ lmin = 8.0e-07 lmax = 1e-06 wmin = 1.5e-05 wmax = 2.0e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.05218230960929+0*(0.0/sqrt(l*w*mult))} lvth0 = 9.14550562624264e-08 wvth0 = -1.8451970633512e-08 pvth0 = 1.24476993893819e-14
+ k1 = 0.589711379999999 lk1 = -9.02707894799971e-9
+ k2 = 0.0185336862874466 lk2 = 1.02256635104885e-08 wk2 = -1.25974239510879e-07 pk2 = 8.49822219740384e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 12212.779 lvsat = 0.0312024228865999
+ ua = -7.09493231346775e-10 lua = 2.06191033386653e-15 wua = 1.78269760282085e-16 pua = -1.20260780286348e-22
+ ub = -6.73962450813236e-21 lub = -1.77838305306815e-25 wub = 7.93645616905948e-23 pub = -5.35393333164753e-29
+ uc = 5.75692682e-12 luc = -5.547051512772e-18 wuc = 2.46519032881566e-32 puc = -1.17549435082229e-38
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0118325541559233 lu0 = 4.40813716641409e-09 wu0 = 1.70585832511132e-07 pu0 = -1.1507720261201e-13
+ a0 = 0.887094242018696 la0 = -2.94019296658117e-08 wa0 = -1.31378030910695e-06 pa0 = 8.86276196523565e-13
+ keta = -0.150384786 lketa = 5.74724026356001e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.962304439039761 lags = -1.62703022576224e-07 wags = -2.08929027487595e-06 pags = 1.40943521943133e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.094399689596+0*(0.009/sqrt(l*w*mult))} lvoff = 1.45567607088616e-8
+ nfactor = {-0.121660262524916+0*(0.02/sqrt(l*w*mult))} lnfactor = 1.33694269509931e-06 wnfactor = 1.71207927521062e-05 pnfactor = -1.15496867905708e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -1.1865e-05 lcit = 1.4750129e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -0.00024405129662779 leta0 = 2.03039284305792e-10 weta0 = 3.55279514569496e-09 peta0 = -2.39671560528582e-15
+ etab = 0.000717673209999999 letab = -6.27676989466e-10
+ dsub = 1.45264382 ldsub = -7.94559948972001e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.98189989655 lpclm = -6.81138389522631e-7
+ pdiblc1 = 0.20581194057 lpdiblc1 = 1.69422666217479e-7
+ pdiblc2 = -0.0319025077049 lpdiblc2 = 2.92192423773255e-08 wpdiblc2 = 2.11758236813575e-22 ppdiblc2 = 5.04870979341448e-29
+ pdiblcb = -0.025
+ drout = 0.33949907438 ldrout = 6.22630675332523e-8
+ pscbe1 = -39572648.0999994 lpscbe1 = 296.53570840826
+ pscbe2 = 1.8099436842e-08 lpscbe2 = -3.10034141461319e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.00023839585627 lalpha0 = -1.49191625283142e-10
+ alpha1 = 0.0
+ beta0 = 66.364220735 lbeta0 = -1.4178399249831e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 4.20616376540937e-08 lagidl = -2.07113247614516e-14 wagidl = -6.59947909687038e-13 pagidl = 4.45200859874876e-19
+ bgidl = 104724742.683838 lbgidl = 1148.55726858548 wbgidl = 17819.3316403754 pbgidl = -0.0120209211245972
+ cgidl = 2177.25520345037 lcgidl = -0.00111798436024762 wcgidl = -0.034921672421848 pcgidl = 2.35581602157787e-8
+ egidl = 1.78393816687 legidl = -8.78937147408501e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.545808072092001 lkt1 = -6.59029745667375e-08 wkt1 = -1.31799790239464e-06 pkt1 = 8.8912138495542e-13
+ kt2 = -0.019032
+ at = 19682.7888368 lat = 0.00358699065069468 wat = 0.52719916095785 pat = -3.55648553982166e-7
+ ute = -2.0356083 lute = 3.74948279179999e-7
+ ua1 = -2.73723400000006e-11 lua1 = 3.91114420564e-16
+ ub1 = -4.5332815e-18 lub1 = 6.35730559899996e-25
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.41e-6
+ sbref = 2.41e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.14 pmos
* DC IV MOS Parameters
+ lmin = 6e-07 lmax = 8.0e-07 wmin = 1.5e-05 wmax = 2.0e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.866730167+0*(0.0/sqrt(l*w*mult))} lvth0 = -3.36509591418e-8
+ k1 = 0.593154569999999 lk1 = -1.1349854922e-8
+ k2 = 0.0156090654 lk2 = 1.219861276116e-8
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 59706.6044000001 lvsat = -0.000836911728239964
+ ua = -1.7341739129e-09 lua = 2.75315992164234e-15
+ ub = 2.4292250742e-18 lub = -1.82114009105532e-24 wub = -1.17549435082229e-38
+ uc = 2.4254276e-12 luc = -3.29962213896e-18
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.00753591610000001 lu0 = 7.30664919894002e-9
+ a0 = 0.932568689999998 la0 = -6.00789922740004e-8
+ keta = 0.0100696950000001 lketa = -5.0770190247e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = -0.533912240000001 lags = 8.46644749104e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {0.00559779755700018+0*(0.009/sqrt(l*w*mult))} lvoff = -5.29015441245522e-8
+ nfactor = {1.7678603+0*(0.02/sqrt(l*w*mult))} lnfactor = 6.2272123620001e-8
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -0.056074191601999 leta0 = 3.78660519343092e-08 weta0 = 1.96868985787621e-22 peta0 = -5.67979851759128e-29
+ etab = -0.00071767321 letab = 3.40607705466e-10
+ dsub = 0.19513736522 ldsub = 5.37539054225879e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.272763882949999 lpclm = 4.71844765251929e-7
+ pdiblc1 = 0.19544523505 lpdiblc1 = 1.7641604576127e-7
+ pdiblc2 = 0.0256746597612 lpdiblc2 = -9.62231479530552e-9
+ pdiblcb = -0.025
+ drout = -0.65870811482 ldrout = 7.35653637367571e-7
+ pscbe1 = 430031833.719999 lpscbe1 = -20.2594750275121
+ pscbe2 = 1.0746893781e-08 lpscbe2 = 1.85968413433741e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -0.000112188837415 lalpha0 = 8.7312809076759e-11 walpha0 = 4.13590306276514e-25 palpha0 = -3.94430452610506e-31
+ alpha1 = 0.0
+ beta0 = 27.750617018 lbeta0 = 1.18703378176572e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 2.28427097e-08 lagidl = -7.74623596362001e-15
+ bgidl = 2044837300 lbgidl = -160.24266258
+ cgidl = 1208.17 lcgidl = -0.000464239482
+ egidl = -0.1972262296 legidl = 4.57556354450159e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.702872459999998 lkt1 = 4.00526615159997e-8
+ kt2 = -0.019032
+ at = 41611.0 lat = -0.0112057806
+ ute = -1.6043825 lute = 8.40433545000009e-8
+ ua1 = 5.53349199999999e-10 lua1 = -6.40330320000131e-19
+ ub1 = -4.2831041e-18 lub1 = 4.66960885859997e-25
+ uc1 = -2.69861592e-10 luc1 = 1.083823099632e-16 wuc1 = 3.15544362088405e-30
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.02e-6
+ sbref = 2.01e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.15 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 6e-07 wmin = 1.5e-05 wmax = 2.0e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.672843265278082+0*(0.0/sqrt(l*w*mult))} lvth0 = -1.25669682699022e-07 wvth0 = -3.46858626146582e-06 pvth0 = 1.64619103969169e-12
+ k1 = 0.4613552 lk1 = 5.12021260800005e-8
+ k2 = 0.0644220228797809 lk2 = -1.09680168587441e-08 wk2 = -5.46221610994454e-07 pk2 = 2.59236776577968e-13
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 47542.9565590052 lvsat = 0.00493595553709614 wvsat = -0.179876037750386 pvsat = 8.53691675163341e-8
+ ua = 1.12102280798156e-08 lua = -3.39025326410048e-15 wua = 3.19039484982239e-17 pua = -1.51416139573701e-23
+ ub = -5.63972439467252e-18 lub = 2.00838332687158e-24 wub = -3.3382969396205e-23 pub = 1.58435572754389e-29
+ uc = -1.70064299999999e-12 luc = -1.3413890322e-18
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0401829011397698 lu0 = -8.18760990093471e-09 wu0 = -8.33896820753414e-08 pu0 = 3.95767431129575e-14
+ a0 = 0.230369639999999 la0 = 2.73184676856001e-7
+ keta = -0.13824211 lketa = 1.9618592406e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 1.25
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.12209155362+0*(0.009/sqrt(l*w*mult))} lvoff = 7.69982194405203e-9
+ nfactor = {-3.32740509415592+0*(0.02/sqrt(l*w*mult))} lnfactor = 2.4804850796864e-06 wnfactor = 9.31941228977392e-05 pnfactor = -4.4229930727267e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 2.873e-05 lcit = -8.88925800000001e-12
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -0.313643296349145 leta0 = 1.60108349047305e-07 weta0 = 2.53081927078373e-06 peta0 = -1.20112682591396e-12
+ etab = 0.0144232238 letab = -6.84526201548001e-9
+ dsub = 0.416017169560001 ldsub = -5.10756497171759e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.006081441 lpclm = 1.23812252201402e-7
+ pdiblc1 = 1.59030588952 lpdiblc1 = -4.85584820850193e-7
+ pdiblc2 = 0.00764468105400001 lpdiblc2 = -1.0652869008684e-9
+ pdiblcb = -0.025
+ drout = 0.860389016439999 ldrout = 1.46901388715754e-8
+ pscbe1 = 479887042.4 lpscbe1 = -43.9207570670401
+ pscbe2 = 1.5334308648e-08 lpscbe2 = -3.17502961540804e-16
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -2.31891527040001e-05 lalpha0 = 4.50735587129184e-11
+ alpha1 = 0.0
+ beta0 = 45.559628338 lbeta0 = 3.41818104518518e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -2.3554226735904e-08 lagidl = 1.42737500688601e-14 wagidl = 4.96770377919715e-14 pagidl = -2.35767221360698e-20
+ bgidl = 2110793275.816 lbgidl = -191.545368702275 wbgidl = -1129.02358618117 pbgidl = 0.000535834594001583
+ cgidl = -8492.23037708105 lcgidl = 0.00413957053696266 wcgidl = 0.126297094444571 pcgidl = -5.99406010233935e-8
+ egidl = 1.1474310464 legidl = -1.80617988739439e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.524531848367999 lkt1 = -4.45877927645482e-08 wkt1 = -2.25804717236236e-06 pkt1 = 1.07166918800318e-12
+ kt2 = -0.019032
+ at = 18000.0
+ ute = -1.6329554 lute = 9.76040528399988e-8
+ ua1 = 5.52e-10
+ ub1 = -7.56664320000001e-18 lub1 = 2.02532854272e-24
+ uc1 = -4.1496e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 1.81e-6
+ sbref = 1.81e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.16 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 1.0e-05 wmax = 1.5e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.964555+0*(0.0/sqrt(l*w*mult))}
+ k1 = 0.59521
+ k2 = 0.02039548
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200000.0
+ ua = 2.7054732e-9
+ ub = -5.157e-20
+ uc = -3.9972e-11
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0209529
+ a0 = 0.8941253
+ keta = -0.0079259
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.1386898
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.093204657+0*(0.009/sqrt(l*w*mult))}
+ nfactor = {1.79934+0*(0.02/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.080000000000001
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.08353125
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0029407877
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 333712830.0
+ pscbe2 = 1.5000958e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 5.0667189e-5
+ alpha1 = 0.0
+ beta0 = 38.266046
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 7.3657e-9
+ bgidl = 1704700000.0
+ cgidl = 700.0
+ egidl = 0.69350825
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.57573
+ kt2 = -0.019032
+ at = 430000.0
+ ute = -1.3864
+ ua1 = 7.0656e-10
+ ub1 = -3.145e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.17 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 1.0e-05 wmax = 1.5e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.964555+0*(0.0/sqrt(l*w*mult))}
+ k1 = 0.59521
+ k2 = 0.02039548
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200000.0
+ ua = 2.7054732e-9
+ ub = -5.157e-20
+ uc = -3.9972e-11
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0209529
+ a0 = 0.8941253
+ keta = -0.0079259
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.1386898
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.093204657+0*(0.009/sqrt(l*w*mult))}
+ nfactor = {1.79934+0*(0.02/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.080000000000001
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.08353125
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0029407877
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 333712830.0
+ pscbe2 = 1.5000958e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 5.0667189e-5
+ alpha1 = 0.0
+ beta0 = 38.266046
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 7.3657e-9
+ bgidl = 1704700000.0
+ cgidl = 700.0
+ egidl = 0.69350825
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.57573
+ kt2 = -0.019032
+ at = 430000.0
+ ute = -1.3864
+ ua1 = 7.0656e-10
+ ub1 = -3.145e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.18 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 1.0e-05 wmax = 1.5e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.9708996575+0*(0.0/sqrt(l*w*mult))} lvth0 = 4.99616399494966e-8
+ k1 = 0.604073147499999 lk1 = -6.9793741303501e-8
+ k2 = 0.017946422832 lk2 = 1.92853455751327e-8
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 296855.3135 lvsat = -0.7626968516871
+ ua = 2.452507249685e-09 lua = 1.99200567235051e-15
+ ub = 2.05160996e-19 lub = -2.0216539011016e-24 pub = 2.80259692864963e-45
+ uc = -5.147278145e-11 luc = 9.05640536061701e-17
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.020337710385 lu0 = 4.84437214227894e-9
+ a0 = 0.913768069025 la0 = -1.54678948964266e-7
+ keta = -0.00498304443500001 lketa = -2.3173810432149e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.113393989575 lags = 1.99194388772705e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0947625464815+0*(0.009/sqrt(l*w*mult))} lvoff = 1.22677565110203e-8
+ nfactor = {1.8039023415+0*(0.02/sqrt(l*w*mult))} lnfactor = -3.59266143759023e-8
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.080000000000001
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.641832441643 lpclm = 5.71194892621197e-06 wpclm = -8.470329472543e-22 ppclm = 6.46234853557053e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 0.004539823205605 lpdiblc2 = -1.25917649924371e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 560098762.7795 lpscbe1 = -1782.69866626545
+ pscbe2 = -1.50486592213e-08 lpscbe2 = 2.36628715770849e-13 ppscbe2 = 3.85185988877447e-34
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 7.7909598465e-05 lalpha0 = -2.14523077573089e-10
+ alpha1 = 0.0
+ beta0 = 39.13253926505 lbeta0 = -6.82328786496286e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 6.546125235e-09 lagidl = 6.45382344446901e-15
+ bgidl = 1480360660.0 lbgidl = 1766.582566764
+ cgidl = 930.5387 lcgidl = -0.00181540004702
+ egidl = 1.2047468705955 legidl = -4.02579964174133e-06 pegidl = -2.58493941422821e-26
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.5851549645 lkt1 = 7.42178254517013e-8
+ kt2 = -0.019032
+ at = 670893.5685 lat = -1.8969404945101
+ ute = -1.222020095 lute = -1.294425999913e-6
+ ua1 = 1.3695660536e-09 lua1 = -5.22090746967856e-15
+ ub1 = -2.61514845e-18 lub1 = -4.17236901562999e-24
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.19 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 1.0e-05 wmax = 1.5e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.9431553561+0*(0.0/sqrt(l*w*mult))} lvth0 = -5.75364302549401e-8
+ k1 = 0.602294036 lk1 = -6.29003958856006e-8
+ k2 = 0.023211373013 lk2 = -1.11423039616984e-9
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 84825.74 lvsat = 0.0588329337960001
+ ua = 3.31328698619e-09 lua = -1.34317149471177e-15
+ ub = -1.239166271e-18 lub = 3.5745365276166e-24 pub = -5.60519385729927e-45
+ uc = -5.44361927e-11 luc = 1.0204608683542e-16
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.02075923934 lu0 = 3.21111605323606e-9
+ a0 = 0.825992817277999 la0 = 1.85415041454661e-7
+ keta = -0.0051939812 lketa = -2.235651484248e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.13791869307 lags = 1.04170972610978e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0645862731911+0*(0.009/sqrt(l*w*mult))} lvoff = -1.04653231979964e-7
+ nfactor = {2.231805466+0*(0.02/sqrt(l*w*mult))} lnfactor = -1.6938800605636e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.020200260000001 leta0 = 2.31700072604e-7
+ etab = -0.1214502716 letab = 1.9934922234136e-7
+ dsub = 0.810118505 ldsub = -9.69109159473e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.044838468325 lpclm = -8.23226181550045e-7
+ pdiblc1 = 0.57808555402 lpdiblc1 = -7.28756287605892e-7
+ pdiblc2 = -0.0010893622944 lpdiblc2 = 9.21907714588223e-09 ppdiblc2 = 2.52435489670724e-29
+ pdiblcb = 0.16246 lpdiblcb = -7.26332516e-07 ppdiblcb = -1.61558713389263e-27
+ drout = 0.147588 ldrout = 1.5979315352e-6
+ pscbe1 = -151521249.434 lpscbe1 = 974.544233056976 ppscbe1 = -1.73472347597681e-18
+ pscbe2 = 7.55293005675e-08 lpscbe2 = -1.14324647226836e-13
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 4.36726325897e-05 lalpha0 = -8.18685295926516e-11
+ alpha1 = -9.37299999999999e-11 lalpha1 = 3.63166258e-16
+ beta0 = 69.5879243857 lbeta0 = -0.000124825723053433
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 9.17928106e-09 lagidl = -3.74860211507602e-15
+ bgidl = 2607594260.0 lbgidl = -2600.996739796
+ cgidl = 455.860685 lcgidl = 2.37873898990002e-5
+ egidl = -1.553543708466 legidl = 6.66147303589036e-06 wegidl = -1.6940658945086e-21 pegidl = -9.69352280335579e-27
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.5669373 lkt1 = 3.63166258000002e-9
+ kt2 = -0.019032
+ at = 209907.023 lat = -0.1108020253158
+ ute = -1.70241253 lute = 5.66902528737998e-7
+ ua1 = -4.749579392e-10 lua1 = 1.92588519282432e-15 wua1 = 5.91645678915759e-31 pua1 = -2.25694915357879e-36
+ ub1 = -3.71946289e-18 lub1 = 1.06407713594007e-25
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.20 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 1.0e-05 wmax = 1.5e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.958701221743304+0*(0.0/sqrt(l*w*mult))} lvth0 = -2.83941505200018e-08 wvth0 = -5.69185171297215e-07 pvth0 = 1.06699452211375e-12
+ k1 = 0.55942551 lk1 = 1.74609429539999e-8
+ k2 = 0.0186737554365172 lk2 = 7.39198751270494e-09 wk2 = -1.5580618679732e-08 pk2 = 2.92074277770254e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 175963.5466 lvsat = -0.11201399845636
+ ua = 3.42372221601093e-09 lua = -1.55019337653409e-15 wua = 6.55553408426568e-18 pua = -1.22890041943799e-23
+ ub = -2.28435241915574e-19 lub = 1.67982014049494e-24 wub = 9.14975067474612e-24 pub = -1.71521226148791e-29
+ uc = 5.12043316e-13 luc = -9.598764001736e-19
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0218668211377404 lu0 = 1.13484321519179e-09 wu0 = 4.86419572560459e-08 pu0 = -9.1184213072184e-14
+ a0 = 0.989848854673976 la0 = -1.21749486247835e-07 wa0 = 2.25481847209484e-07 pa0 = -4.2268827077889e-13
+ keta = 0.0419609792 lketa = -1.1075320360832e-07 pketa = 2.01948391736579e-28
+ a1 = 0.0
+ a2 = 0.5
+ ags = -0.313790559479661 lags = 9.50945137440573e-07 wags = 3.8139368322653e-07 pags = -7.14960598576452e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1577214518922+0*(0.009/sqrt(l*w*mult))} lvoff = 6.99379740131182e-8
+ nfactor = {1.23095735709116+0*(0.02/sqrt(l*w*mult))} lnfactor = 1.82309804396918e-07 wnfactor = -2.99753248679908e-06 pnfactor = 5.61917439975356e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.4373e-05 lcit = -8.19762580000001e-12
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.269530642722601 leta0 = -2.35694662847786e-7
+ etab = -0.0283214568 letab = 2.476994611728e-8
+ dsub = 0.0736166540000001 ldsub = 4.115372104116e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.0832187031859539 lpclm = 9.79426230179612e-07 wpclm = -3.30153811658551e-10 ppclm = 6.18906335329684e-16
+ pdiblc1 = 0.00549710251999991 lpdiblc1 = 3.44618023576008e-7
+ pdiblc2 = 0.00585964945018 lpdiblc2 = -3.80754027050743e-9
+ pdiblcb = -0.39992 lpdiblcb = 3.27905032e-7
+ drout = 1.515411042014 ldrout = -9.66189539359445e-7
+ pscbe1 = 428577028.488 lpscbe1 = -112.907998735605
+ pscbe2 = 1.45331535696e-08 lpscbe2 = 1.87299354278452e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -5.93092031506e-05 lalpha0 = 1.11181219686115e-10 walpha0 = 4.52253956963206e-26 palpha0 = -1.91361452517254e-31
+ alpha1 = 1.8746e-10 lalpha1 = -1.63952516e-16
+ beta0 = -38.239948205 lbeta0 = 7.7308406905093e-05 wbeta0 = -2.71050543121376e-20
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 6.15911672e-09 lagidl = 1.912997956688e-15
+ bgidl = 810087519.999999 lbgidl = 768.609395008
+ cgidl = 556.49103 lcgidl = -0.000164854254838
+ egidl = 3.067904826664 legidl = -2.00189438806434e-6
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.478686475497216 lkt1 = -1.61803333032919e-07 wkt1 = -2.95817815244957e-07 pkt1 = 5.54540076458189e-13
+ kt2 = -0.019032
+ at = 251716.309990624 lat = -0.189177714708424 wat = 0.0475421488786534 pat = -8.91225122879235e-8
+ ute = -0.962470120905648 lute = -8.20193511350274e-07 wute = -3.85883775065069e-06 pute = 7.23377724736976e-12
+ ua1 = 9.01186308801705e-10 lua1 = -6.53834814479677e-16 wua1 = -3.50174338796213e-15 pua1 = 6.56436815507381e-21
+ ub1 = -3.15856725943304e-18 lub1 = -9.45047235466823e-25 wub1 = -5.69185171297205e-24 pub1 = 1.06699452211375e-29
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.81e-6
+ sbref = 2.81e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.21 pmos
* DC IV MOS Parameters
+ lmin = 8.0e-07 lmax = 1e-06 wmin = 1.0e-05 wmax = 1.5e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.24263554628348+0*(0.0/sqrt(l*w*mult))} lvth0 = 2.19934809722836e-07 wvth0 = 2.84592585648606e-06 pvth0 = -1.91986158278549e-12
+ k1 = 0.589711380000001 lk1 = -9.02707894799971e-9
+ k2 = 0.0049778286874142 lk2 = 1.93704450474703e-08 wk2 = 7.79030933986593e-08 pk2 = -5.25534268067355e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 12212.779 lvsat = 0.0312024228866
+ ua = -6.9546063205464e-10 lua = 2.05244394238406e-15 wua = -3.27776704213536e-17 pua = 2.2111816466258e-23
+ ub = 8.31207766957787e-18 lub = -5.78971245189723e-24 wub = -4.57487533737306e-23 pub = 3.08621090259186e-29
+ uc = 5.75692682e-12 luc = -5.547051512772e-18
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0393459339112979 lu0 = -1.41523888165615e-08 wu0 = -2.4320978628023e-07 pu0 = 1.64069321824643e-13
+ a0 = 0.87470238025012 la0 = -2.10423797167305e-08 wa0 = -1.1274092360474e-06 pa0 = 7.60550270637573e-13
+ keta = -0.150384786 lketa = 5.74724026356e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.950181810598304 lags = -1.54525097429615e-07 wags = -1.90696841613265e-06 pags = 1.28644089352307e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0943996895960002+0*(0.009/sqrt(l*w*mult))} lvoff = 1.45567607088615e-8
+ nfactor = {0.0201721345442181+0*(0.02/sqrt(l*w*mult))} lnfactor = 1.24126256003647e-06 wnfactor = 1.49876624339954e-05 pnfactor = -1.01106770779733e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -1.1865e-05 lcit = 1.4750129e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -7.82501099898989e-06 leta0 = 4.36810320206e-11
+ etab = 0.00071767321 letab = -6.27676989466e-10
+ dsub = 1.45264382 ldsub = -7.94559948972e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.98179013648023 lpclm = -6.81064345379564e-07 wpclm = 1.65076905828598e-09 ppclm = -1.11360880671717e-15
+ pdiblc1 = 0.20581194057 lpdiblc1 = 1.69422666217478e-7
+ pdiblc2 = -0.0319025077049 lpdiblc2 = 2.92192423773255e-08 wpdiblc2 = -1.05879118406788e-22 ppdiblc2 = -2.52435489670724e-29
+ pdiblcb = -0.025
+ drout = 0.33949907438 ldrout = 6.22630675332523e-8
+ pscbe1 = -39572648.0999999 lpscbe1 = 296.535708408259
+ pscbe2 = 1.8099436842e-08 lpscbe2 = -3.10034141461319e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.00023839585627 lalpha0 = -1.49191625283142e-10
+ alpha1 = 0.0
+ beta0 = 66.3642207350001 lbeta0 = -1.4178399249831e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -1.8184728e-09 lagidl = 8.89019775088e-15
+ bgidl = 1289536800 lbgidl = 349.283054719999
+ cgidl = -144.695999999999 lcgidl = 0.0004484039216
+ egidl = 1.78393816687 legidl = -8.78937147408503e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.73178712251392 lkt1 = 5.95584928478902e-08 wkt1 = 1.47908907622477e-06 pkt1 = -9.97793490821222e-13
+ kt2 = -0.019032
+ at = 70541.85004688 lat = -0.0307225320416252 wat = -0.237710744393266 pat = 1.60359668167697e-7
+ ute = -3.31848399547176 lute = 1.24037622334525e-06 wute = 1.92941887532534e-05 pute = -1.30158597329447e-11
+ ua1 = -1.19153154400853e-09 lua1 = 1.17645621958815e-15 wua1 = 1.75087169398106e-14 pua1 = -1.18113804475962e-20
+ ub1 = -6.4255451028348e-18 lub1 = 1.91225158637235e-24 wub1 = 2.84592585648604e-23 pub1 = -1.91986158278548e-29
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.41e-6
+ sbref = 2.41e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.22 pmos
* DC IV MOS Parameters
+ lmin = 6e-07 lmax = 8.0e-07 wmin = 1.0e-05 wmax = 1.5e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.866730167+0*(0.0/sqrt(l*w*mult))} lvth0 = -3.36509591418e-8
+ k1 = 0.593154570000001 lk1 = -1.1349854922e-8
+ k2 = 0.0156090654 lk2 = 1.219861276116e-8
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 59706.6044 lvsat = -0.00083691172824002
+ ua = -1.7341739129e-09 lua = 2.75315992164234e-15
+ ub = 2.4292250742e-18 lub = -1.82114009105532e-24 wub = 5.87747175411144e-39 pub = -2.80259692864963e-45
+ uc = 2.4254276e-12 luc = -3.29962213896e-18
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.00753591610000001 lu0 = 7.30664919894001e-9
+ a0 = 0.932568689999998 la0 = -6.00789922739996e-8
+ keta = 0.010069695 lketa = -5.0770190247e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = -0.53391224 lags = 8.46644749104e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {0.00559779755700007+0*(0.009/sqrt(l*w*mult))} lvoff = -5.29015441245523e-8
+ nfactor = {1.7678603+0*(0.02/sqrt(l*w*mult))} lnfactor = 6.22721236199993e-8
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -0.056074191601999 leta0 = 3.78660519343092e-08 weta0 = 9.0989867380833e-24 peta0 = 4.77260847658712e-29
+ etab = -0.00071767321 letab = 3.40607705466e-10
+ dsub = 0.19513736522 ldsub = 5.37539054225877e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.272763882950001 lpclm = 4.7184476525193e-7
+ pdiblc1 = 0.195445235049999 lpdiblc1 = 1.7641604576127e-7
+ pdiblc2 = 0.0256746597612 lpdiblc2 = -9.62231479530552e-9
+ pdiblcb = -0.025
+ drout = -0.65870811482 ldrout = 7.35653637367572e-7
+ pscbe1 = 430031833.72 lpscbe1 = -20.2594750275121
+ pscbe2 = 1.0746893781e-08 lpscbe2 = 1.85968413433741e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -0.000112188837415 lalpha0 = 8.7312809076759e-11 walpha0 = 2.06795153138257e-25 palpha0 = -9.86076131526265e-32
+ alpha1 = 0.0
+ beta0 = 27.750617018 lbeta0 = 1.18703378176572e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 2.28427097e-08 lagidl = -7.74623596362001e-15
+ bgidl = 2044837300.0 lbgidl = -160.24266258
+ cgidl = 1208.17 lcgidl = -0.000464239482 wcgidl = 6.93889390390723e-18
+ egidl = -0.197226229600001 legidl = 4.5755635445016e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.70287246 lkt1 = 4.00526615160001e-8
+ kt2 = -0.019032
+ at = 41611.0 lat = -0.0112057806
+ ute = -1.6043825 lute = 8.40433545e-8
+ ua1 = 5.53349200000001e-10 lua1 = -6.40330319999736e-19
+ ub1 = -4.2831041e-18 lub1 = 4.66960885859997e-25
+ uc1 = -2.69861592e-10 luc1 = 1.083823099632e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.02e-6
+ sbref = 2.01e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.23 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 6e-07 wmin = 1.0e-05 wmax = 1.5e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.936303203187368+0*(0.0/sqrt(l*w*mult))} lvth0 = -6.31596167274917e-10 wvth0 = 4.93797458862491e-07 pvth0 = -2.34356273976135e-13
+ k1 = 0.4613552 lk1 = 5.12021260800001e-8
+ k2 = 0.0165801831699776 lk2 = 1.17377202675286e-08 wk2 = 1.73309898505689e-07 pk2 = -8.22528778307995e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 39062.5430944962 lvsat = 0.00896075976735206 wvsat = -0.0523323492485179 pvsat = 2.48369329533469e-8
+ ua = 1.12059934479471e-08 lua = -3.38824350781569e-15 wua = 9.55919479355897e-17 pua = -4.53679384902738e-23
+ ub = -1.0140432494792e-17 lub = 4.1444193911883e-24 wub = 3.43067622851402e-23 pub = -1.62819893805275e-29
+ uc = -1.70064299999999e-12 luc = -1.3413890322e-18
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0279596795165948 lu0 = -2.38646891857587e-09 wu0 = 1.004450776e-07 pu0 = -4.767123382896e-14
+ a0 = 0.230369639999999 la0 = 2.73184676856e-7
+ keta = -0.13824211 lketa = 1.9618592406e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 1.25
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.12209155362+0*(0.009/sqrt(l*w*mult))} lvoff = 7.69982194405203e-9
+ nfactor = {6.49889904330542+0*(0.02/sqrt(l*w*mult))} lnfactor = -2.18307886395275e-06 wnfactor = -5.45914867636355e-05 pnfactor = 2.59091196180214e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 2.873e-05 lcit = -8.88925800000001e-12
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -0.181495734228849 leta0 = 9.73911160650121e-08 weta0 = 5.43346894597139e-07 peta0 = -2.57872436175802e-13
+ etab = -0.0116421222850369 letab = 5.52535123647852e-09 wetab = 3.92017487788354e-07 petab = -1.86051499704353e-13
+ dsub = 0.41601716956 ldsub = -5.10756497171763e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.201999400053921 lpclm = 5.05429588834408e-07 wpclm = 1.20932298630927e-05 ppclm = -5.73944689302379e-12
+ pdiblc1 = 1.59030588952 lpdiblc1 = -4.85584820850192e-7
+ pdiblc2 = 0.007644681054 lpdiblc2 = -1.0652869008684e-9
+ pdiblcb = -0.025
+ drout = 0.860389016440001 ldrout = 1.46901388715754e-8
+ pscbe1 = 479887042.4 lpscbe1 = -43.9207570670401
+ pscbe2 = 1.5334308648e-08 lpscbe2 = -3.17502961540804e-16
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -2.31891527040001e-05 lalpha0 = 4.50735587129185e-11
+ alpha1 = 0.0
+ beta0 = 45.559628338 lbeta0 = 3.41818104518518e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -6.66457433266176e-08 lagidl = 3.47249838428127e-14 wagidl = 6.97764656646919e-13 pagidl = -3.31159106044628e-19
+ bgidl = 1567115115.33264 lbgidl = 66.4842862631303 wbgidl = 7047.78503714383 pbgidl = -0.00334487877862846
+ cgidl = -487.342031519039 lcgidl = 0.000340450528158936 wcgidl = 0.00590520672454105 pcgidl = -2.80261111146718e-9
+ egidl = 1.1474310464 legidl = -1.8061798873944e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.674670000000001 lkt1 = 2.66677739999999e-8
+ kt2 = -0.019032
+ at = 18000.0
+ ute = -1.6329554 lute = 9.76040528399996e-8
+ ua1 = 5.52e-10
+ ub1 = -7.56664320000001e-18 lub1 = 2.02532854272e-24
+ uc1 = -4.1496e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 1.81e-6
+ sbref = 1.81e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.24 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 7e-06 wmax = 1.0e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.964555+0*(0.0/sqrt(l*w*mult))}
+ k1 = 0.59521
+ k2 = 0.02039548
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200000.0
+ ua = 2.7054732e-9
+ ub = -5.157e-20
+ uc = -3.9972e-11
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0209529
+ a0 = 0.8941253
+ keta = -0.0079259
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.1386898
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.093204657+0*(0.009/sqrt(l*w*mult))}
+ nfactor = {1.79934+0*(0.02/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.080000000000001
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.08353125
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0029407877
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 333712830.0
+ pscbe2 = 1.5000958e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 5.0667189e-5
+ alpha1 = 0.0
+ beta0 = 38.266046
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 7.3657e-9
+ bgidl = 1704700000.0
+ cgidl = 700.0
+ egidl = 0.69350825
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.57573
+ kt2 = -0.019032
+ at = 430000.0
+ ute = -1.3864
+ ua1 = 7.0656e-10
+ ub1 = -3.145e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.25 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 7e-06 wmax = 1.0e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.964555+0*(0.0/sqrt(l*w*mult))}
+ k1 = 0.59521
+ k2 = 0.02039548
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200000.0
+ ua = 2.7054732e-9
+ ub = -5.157e-20
+ uc = -3.9972e-11
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0209529
+ a0 = 0.8941253
+ keta = -0.0079259
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.1386898
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.093204657+0*(0.009/sqrt(l*w*mult))}
+ nfactor = {1.79934+0*(0.02/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.080000000000001
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.08353125
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0029407877
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 333712830.0
+ pscbe2 = 1.5000958e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 5.0667189e-5
+ alpha1 = 0.0
+ beta0 = 38.266046
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 7.3657e-9
+ bgidl = 1704700000.0
+ cgidl = 700.0
+ egidl = 0.69350825
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.57573
+ kt2 = -0.019032
+ at = 430000.0
+ ute = -1.3864
+ ua1 = 7.0656e-10
+ ub1 = -3.145e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.26 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 7e-06 wmax = 1.0e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.9708996575+0*(0.0/sqrt(l*w*mult))} lvth0 = 4.99616399494966e-8
+ k1 = 0.6040731475 lk1 = -6.97937413034993e-8
+ k2 = 0.017946422832 lk2 = 1.92853455751329e-8
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 296855.3135 lvsat = -0.7626968516871
+ ua = 2.452507249685e-09 lua = 1.9920056723505e-15
+ ub = 2.05160996e-19 lub = -2.0216539011016e-24 pub = -1.40129846432482e-45
+ uc = -5.147278145e-11 luc = 9.05640536061702e-17
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.020337710385 lu0 = 4.84437214227894e-9
+ a0 = 0.913768069025 la0 = -1.54678948964262e-7
+ keta = -0.00498304443499999 lketa = -2.3173810432149e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.113393989575 lags = 1.99194388772705e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0947625464815+0*(0.009/sqrt(l*w*mult))} lvoff = 1.22677565110203e-8
+ nfactor = {1.8039023415+0*(0.02/sqrt(l*w*mult))} lnfactor = -3.59266143759023e-8
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.080000000000001
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.641832441643 lpclm = 5.71194892621197e-06 wpclm = 8.470329472543e-22 ppclm = -6.46234853557053e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 0.004539823205605 lpdiblc2 = -1.25917649924371e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 560098762.7795 lpscbe1 = -1782.69866626545
+ pscbe2 = -1.50486592213e-08 lpscbe2 = 2.36628715770849e-13 ppscbe2 = -3.85185988877447e-34
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 7.7909598465e-05 lalpha0 = -2.14523077573089e-10
+ alpha1 = 0.0
+ beta0 = 39.13253926505 lbeta0 = -6.82328786496265e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 6.546125235e-09 lagidl = 6.45382344446901e-15
+ bgidl = 1480360660.0 lbgidl = 1766.582566764
+ cgidl = 930.5387 lcgidl = -0.00181540004702
+ egidl = 1.2047468705955 legidl = -4.02579964174133e-6
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.5851549645 lkt1 = 7.42178254516979e-8
+ kt2 = -0.019032
+ at = 670893.5685 lat = -1.8969404945101
+ ute = -1.222020095 lute = -1.294425999913e-6
+ ua1 = 1.3695660536e-09 lua1 = -5.22090746967856e-15
+ ub1 = -2.61514845e-18 lub1 = -4.17236901563e-24
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.27 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 7e-06 wmax = 1.0e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.943155356100001+0*(0.0/sqrt(l*w*mult))} lvth0 = -5.75364302549384e-8
+ k1 = 0.602294036 lk1 = -6.29003958855998e-8
+ k2 = 0.023211373013 lk2 = -1.11423039616978e-9
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 84825.7400000001 lvsat = 0.0588329337959999
+ ua = 3.31328698619e-09 lua = -1.34317149471177e-15
+ ub = -1.239166271e-18 lub = 3.5745365276166e-24 pub = -5.60519385729927e-45
+ uc = -5.44361927e-11 luc = 1.0204608683542e-16
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.02075923934 lu0 = 3.21111605323603e-9
+ a0 = 0.825992817278001 la0 = 1.85415041454661e-7
+ keta = -0.0051939812 lketa = -2.235651484248e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.13791869307 lags = 1.04170972610978e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0645862731911+0*(0.009/sqrt(l*w*mult))} lvoff = -1.04653231979964e-7
+ nfactor = {2.231805466+0*(0.02/sqrt(l*w*mult))} lnfactor = -1.6938800605636e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.0202002600000011 leta0 = 2.31700072604e-7
+ etab = -0.1214502716 letab = 1.9934922234136e-7
+ dsub = 0.810118505 ldsub = -9.69109159473001e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.044838468325 lpclm = -8.23226181550045e-7
+ pdiblc1 = 0.57808555402 lpdiblc1 = -7.28756287605892e-7
+ pdiblc2 = -0.0010893622944 lpdiblc2 = 9.21907714588224e-09 ppdiblc2 = 1.26217744835362e-29
+ pdiblcb = 0.16246 lpdiblcb = -7.26332516e-07 wpdiblcb = -2.11758236813575e-22 ppdiblcb = -1.21169035041947e-27
+ drout = 0.147588000000001 ldrout = 1.5979315352e-6
+ pscbe1 = -151521249.434 lpscbe1 = 974.544233056976
+ pscbe2 = 7.55293005675e-08 lpscbe2 = -1.14324647226836e-13
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 4.36726325897e-05 lalpha0 = -8.18685295926516e-11
+ alpha1 = -9.37299999999999e-11 lalpha1 = 3.63166258e-16
+ beta0 = 69.5879243857 lbeta0 = -0.000124825723053433
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 9.17928106000001e-09 lagidl = -3.74860211507601e-15
+ bgidl = 2607594260.0 lbgidl = -2600.996739796
+ cgidl = 455.860685 lcgidl = 2.37873898990002e-5
+ egidl = -1.553543708466 legidl = 6.66147303589036e-06 wegidl = 8.470329472543e-22 pegidl = 1.13091099372484e-26
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.5669373 lkt1 = 3.63166258000002e-9
+ kt2 = -0.019032
+ at = 209907.023 lat = -0.1108020253158
+ ute = -1.70241253 lute = 5.66902528738001e-7
+ ua1 = -4.74957939199999e-10 lua1 = 1.92588519282432e-15 wua1 = -1.97215226305253e-31 pua1 = -1.88079096131566e-36
+ ub1 = -3.71946289e-18 lub1 = 1.06407713594001e-25
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.28 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 7e-06 wmax = 1.0e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.0153941238+0*(0.0/sqrt(l*w*mult))} lvth0 = 7.78823636754802e-8
+ k1 = 0.55942551 lk1 = 1.74609429539999e-8
+ k2 = 0.017121869454 lk2 = 1.03011529755316e-8
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 175963.5466 lvsat = -0.11201399845636
+ ua = 3.42437517092e-09 lua = -1.55141740580663e-15
+ ub = 6.82913023999999e-19 lub = -2.85933187904e-26
+ uc = 5.12043316e-13 luc = -9.598764001736e-19
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.02671173604 lu0 = -7.94743426058401e-9
+ a0 = 1.012307662324 la0 = -1.63850767068571e-7
+ keta = 0.0419609792 lketa = -1.1075320360832e-07 pketa = -1.0097419586829e-28
+ a1 = 0.0
+ a2 = 0.5
+ ags = -0.27580236896 lags = 8.79732475492417e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1577214518922+0*(0.009/sqrt(l*w*mult))} lvoff = 6.99379740131181e-8
+ nfactor = {0.932392277999998+0*(0.02/sqrt(l*w*mult))} lnfactor = 7.41999901661201e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.4373e-05 lcit = -8.1976258e-12
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.269530642722601 leta0 = -2.35694662847786e-7
+ etab = -0.0283214568 letab = 2.476994611728e-8
+ dsub = 0.0736166539999998 ldsub = 4.115372104116e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.0831858186719994 lpclm = 9.7948787548947e-7
+ pdiblc1 = 0.00549710251999991 lpdiblc1 = 3.44618023576008e-7
+ pdiblc2 = 0.00585964945018 lpdiblc2 = -3.80754027050743e-9
+ pdiblcb = -0.39992 lpdiblcb = 3.27905032e-7
+ drout = 1.515411042014 ldrout = -9.66189539359445e-7
+ pscbe1 = 428577028.488 lpscbe1 = -112.907998735605 wpscbe1 = 1.81898940354586e-12
+ pscbe2 = 1.45331535696e-08 lpscbe2 = 1.87299354278452e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -5.93092031506e-05 lalpha0 = 1.11181219686115e-10 walpha0 = -2.36279618331797e-26 palpha0 = -8.09153887377223e-32
+ alpha1 = 1.8746e-10 lalpha1 = -1.63952516e-16
+ beta0 = -38.239948205 lbeta0 = 7.7308406905093e-05 pbeta0 = 2.58493941422821e-26
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 6.15911672e-09 lagidl = 1.912997956688e-15
+ bgidl = 810087519.999999 lbgidl = 768.609395008
+ cgidl = 556.49103 lcgidl = -0.000164854254838
+ egidl = 3.067904826664 legidl = -2.00189438806434e-6
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.508151 lkt1 = -1.065691354e-7
+ kt2 = -0.019032
+ at = 256451.68 lat = -0.198054639328 wat = 8.88178419700125e-16
+ ute = -1.34682432 lute = -9.96831297280004e-8
+ ua1 = 5.524e-10
+ ub1 = -3.72549628e-18 lub1 = 1.17717906487999e-25
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.81e-6
+ sbref = 2.81e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.29 pmos
* DC IV MOS Parameters
+ lmin = 8.0e-07 lmax = 1e-06 wmin = 7e-06 wmax = 1.0e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.959171036000001+0*(0.0/sqrt(l*w*mult))} lvth0 = 2.87096510855984e-8
+ k1 = 0.589711379999999 lk1 = -9.02707894799886e-9
+ k2 = 0.0127372586 lk2 = 1.413593362844e-8
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 12212.779 lvsat = 0.0312024228866
+ ua = -6.98725406600002e-10 lua = 2.05464635929236e-15
+ ub = 3.75533634e-18 lub = -2.715734750964e-24 pub = -5.60519385729927e-45
+ uc = 5.75692682e-12 luc = -5.547051512772e-18 puc = -5.87747175411144e-39
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0151213594 lu0 = 2.18950914875996e-9
+ a0 = 0.762408342000001 la0 = 5.47111784867976e-8
+ keta = -0.150384786 lketa = 5.74724026356e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.760240858 lags = -2.63909308067991e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.094399689596+0*(0.009/sqrt(l*w*mult))} lvoff = 1.45567607088615e-8
+ nfactor = {1.51299753+0*(0.02/sqrt(l*w*mult))} lnfactor = 2.34202548261998e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -1.1865e-05 lcit = 1.4750129e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -7.82501099899e-06 leta0 = 4.36810320206e-11
+ etab = 0.00071767321 letab = -6.27676989466e-10
+ dsub = 1.45264382 ldsub = -7.94559948971999e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.98195455905 lpclm = -6.8117526484513e-7
+ pdiblc1 = 0.205811940570001 lpdiblc1 = 1.69422666217478e-7
+ pdiblc2 = -0.0319025077049 lpdiblc2 = 2.92192423773255e-08 wpdiblc2 = -5.29395592033938e-23 ppdiblc2 = 1.26217744835362e-29
+ pdiblcb = -0.025
+ drout = 0.339499074379999 ldrout = 6.22630675332515e-8
+ pscbe1 = -39572648.0999994 lpscbe1 = 296.53570840826
+ pscbe2 = 1.8099436842e-08 lpscbe2 = -3.10034141461319e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.00023839585627 lalpha0 = -1.49191625283142e-10
+ alpha1 = 0.0
+ beta0 = 66.3642207350001 lbeta0 = -1.41783992498309e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -1.81847280000003e-09 lagidl = 8.89019775088e-15
+ bgidl = 1289536800 lbgidl = 349.283054719999
+ cgidl = -144.696000000001 lcgidl = 0.0004484039216
+ egidl = 1.78393816687 legidl = -8.78937147408501e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.584464499999999 lkt1 = -3.98253483000005e-8
+ kt2 = -0.019032
+ at = 46864.9999999999 lat = -0.0147501290000001
+ ute = -1.396713 lute = -5.60504901999988e-8
+ ua1 = 5.524e-10
+ ub1 = -3.5909e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.41e-6
+ sbref = 2.41e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.30 pmos
* DC IV MOS Parameters
+ lmin = 6e-07 lmax = 8.0e-07 wmin = 7e-06 wmax = 1.0e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.866730166999998+0*(0.0/sqrt(l*w*mult))} lvth0 = -3.36509591418008e-8
+ k1 = 0.59315457 lk1 = -1.1349854922e-8
+ k2 = 0.0156090654 lk2 = 1.219861276116e-8
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 59706.6044 lvsat = -0.000836911728240075
+ ua = -1.73417391290001e-09 lua = 2.75315992164234e-15
+ ub = 2.4292250742e-18 lub = -1.82114009105532e-24 wub = -2.93873587705572e-39 pub = 1.40129846432482e-45
+ uc = 2.42542760000001e-12 luc = -3.29962213896e-18
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.00753591609999998 lu0 = 7.30664919893999e-9
+ a0 = 0.93256869 la0 = -6.00789922739996e-8
+ keta = 0.0100696950000001 lketa = -5.0770190247e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = -0.533912239999999 lags = 8.46644749104e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {0.00559779755700007+0*(0.009/sqrt(l*w*mult))} lvoff = -5.29015441245522e-8
+ nfactor = {1.7678603+0*(0.02/sqrt(l*w*mult))} lnfactor = 6.22721236199993e-8
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -0.056074191601999 leta0 = 3.78660519343092e-08 weta0 = -3.22600438895681e-23 peta0 = 3.1948866661451e-29
+ etab = -0.00071767321 letab = 3.40607705466e-10
+ dsub = 0.19513736522 ldsub = 5.37539054225881e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.272763882949999 lpclm = 4.7184476525193e-7
+ pdiblc1 = 0.195445235049999 lpdiblc1 = 1.7641604576127e-7
+ pdiblc2 = 0.0256746597612 lpdiblc2 = -9.62231479530551e-9
+ pdiblcb = -0.025
+ drout = -0.658708114820001 ldrout = 7.35653637367572e-7
+ pscbe1 = 430031833.72 lpscbe1 = -20.2594750275116
+ pscbe2 = 1.0746893781e-08 lpscbe2 = 1.85968413433739e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -0.000112188837415 lalpha0 = 8.73128090767591e-11 walpha0 = 2.06795153138257e-25 palpha0 = 1.97215226305253e-31
+ alpha1 = 0.0
+ beta0 = 27.750617018 lbeta0 = 1.18703378176572e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 2.28427097e-08 lagidl = -7.74623596362e-15 wagidl = 1.0097419586829e-28
+ bgidl = 2044837300 lbgidl = -160.24266258
+ cgidl = 1208.17 lcgidl = -0.000464239482000001
+ egidl = -0.1972262296 legidl = 4.57556354450161e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.702872459999999 lkt1 = 4.00526615160001e-8
+ kt2 = -0.019032
+ at = 41611.0 lat = -0.0112057806
+ ute = -1.6043825 lute = 8.40433545000009e-8
+ ua1 = 5.533492e-10 lua1 = -6.40330319999736e-19
+ ub1 = -4.2831041e-18 lub1 = 4.66960885860003e-25
+ uc1 = -2.69861592e-10 luc1 = 1.083823099632e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.02e-6
+ sbref = 2.01e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.31 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 6e-07 wmin = 7e-06 wmax = 1.0e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.02/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.839378752414435+0*(0.0/sqrt(l*w*mult))} lvth0 = -4.66319405041099e-08 wvth0 = -4.79304254309809e-07 pvth0 = 2.27477799095439e-13
+ k1 = 0.4613552 lk1 = 5.12021260800001e-8
+ k2 = 0.0357851452517788 lk2 = 2.62304526350585e-09 wk2 = -1.9504002983331e-08 pk2 = 9.25659981588866e-15
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 19030.3862272684 lvsat = 0.0184680214165383 wvsat = 0.148786419138448 pvsat = -7.06140345231069e-8
+ ua = 1.12232294341828e-08 lua = -3.39642370688316e-15 wua = -7.74538377297236e-17 pua = 3.67595913865197e-23
+ ub = -5.63493266588763e-18 lub = 2.00610917239027e-24 wub = -1.09275368750949e-23 pub = 5.18620900092005e-30
+ uc = -1.70064300000001e-12 luc = -1.34138903220001e-18
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0328088272779721 lu0 = -4.68787444612554e-09 wu0 = 5.17606233019156e-08 pu0 = -2.45655918190889e-14
+ a0 = 0.230369639999997 la0 = 2.73184676856001e-7
+ keta = -0.13824211 lketa = 1.9618592406e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 1.25
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.12209155362+0*(0.009/sqrt(l*w*mult))} lvoff = 7.69982194405214e-9
+ nfactor = {0.633211112334216+0*(0.02/sqrt(l*w*mult))} lnfactor = 6.00776628086181e-07 wnfactor = 4.29882346297746e-06 pnfactor = -2.04022161552911e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 2.873e-05 lcit = -8.88925800000001e-12
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.0133660136299926 leta0 = 4.90973053120592e-09 weta0 = -1.41302530210907e-06 peta0 = 6.70621808380962e-13
+ etab = 0.0578654672750616 letab = -2.74629507687442e-08 wetab = -3.05824531846764e-07 petab = 1.45144322814474e-13
+ dsub = 0.41601716956 ldsub = -5.10756497171759e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.34650034642137 lpclm = -5.1235056031158e-07 wpclm = -9.4371221602434e-06 ppclm = 4.47885817725151e-12
+ pdiblc1 = 1.59030588952 lpdiblc1 = -4.85584820850192e-7
+ pdiblc2 = 0.007644681054 lpdiblc2 = -1.0652869008684e-9
+ pdiblcb = -0.025
+ drout = 0.860389016439999 ldrout = 1.46901388715754e-8
+ pscbe1 = 479887042.4 lpscbe1 = -43.9207570670401
+ pscbe2 = 1.5334308648e-08 lpscbe2 = -3.17502961540804e-16
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -2.31891527040003e-05 lalpha0 = 4.50735587129184e-11
+ alpha1 = 0.0
+ beta0 = 45.5596283379999 lbeta0 = 3.41818104518518e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 2.65881088344e-08 lagidl = -9.52380239280623e-15 wagidl = -2.38284199343856e-13 pagidl = 1.13089681008594e-19
+ bgidl = 2269100000.0 lbgidl = -266.677740000001
+ cgidl = -694.513726610559 lcgidl = 0.000438774214649372 wcgidl = 0.0079851682802341 pcgidl = -3.78976086579911e-9
+ egidl = 1.1474310464 legidl = -1.8061798873944e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.674670000000001 lkt1 = 2.66677739999999e-8
+ kt2 = -0.019032
+ at = 18000.0
+ ute = -1.6329554 lute = 9.76040528400005e-8
+ ua1 = 5.52e-10
+ ub1 = -7.5666432e-18 lub1 = 2.02532854272e-24
+ uc1 = -4.1496e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 1.81e-6
+ sbref = 1.81e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.32 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.981471075273999+0*(0.0/sqrt(l*w*mult))} wvth0 = 1.19085719049605e-7
+ k1 = 0.59521
+ k2 = 0.02024960310478 wk2 = 1.02694358346211e-9
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200000.0
+ ua = 2.70605602720842e-09 wua = -4.10298465052088e-18
+ ub = 9.72299769e-20 wub = -1.04752148218071e-24
+ uc = -3.9972e-11
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0222478755822 wu0 = -9.11636392366927e-9
+ a0 = 0.892767301768819 wa0 = 9.56003051587095e-9
+ keta = -0.0079259
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.1452740414842 wags = -4.63517168635051e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.093204657+0*(0.009/sqrt(l*w*mult))}
+ nfactor = {1.77182271384+0*(0.02/sqrt(l*w*mult))} wnfactor = 1.93716081040028e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.080000000000001
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.08353125
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0029407877
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 333712830.0
+ pscbe2 = 1.5000958e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 5.0667189e-5
+ alpha1 = 0.0
+ beta0 = 38.266046
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -1.27942399694e-08 wagidl = 1.41921864756822e-13
+ bgidl = 1704700000.0
+ cgidl = -55.9694000000009 wcgidl = 0.0053218703582424
+ egidl = 0.69350825
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.575049627539999 wkt1 = -4.78968332241747e-9
+ kt2 = -0.019032
+ at = 382625.9176 wat = 0.33350387578319
+ ute = -1.0091712694 wute = -2.65561330876296e-6
+ ua1 = 2.431339464672e-09 wua1 = -1.21420955762801e-14
+ ub1 = -1.8404488054e-18 wub1 = -9.1837742815403e-24
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.33 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.981471075274+0*(0.0/sqrt(l*w*mult))} wvth0 = 1.19085719049609e-7
+ k1 = 0.59521
+ k2 = 0.02024960310478 wk2 = 1.02694358346221e-9
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200000.0
+ ua = 2.70605602720842e-09 wua = -4.10298465052088e-18
+ ub = 9.72299769000001e-20 wub = -1.04752148218071e-24
+ uc = -3.9972e-11
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0222478755822 wu0 = -9.11636392366932e-9
+ a0 = 0.89276730176882 wa0 = 9.56003051587095e-9
+ keta = -0.0079259
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.1452740414842 wags = -4.63517168635059e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.093204657+0*(0.009/sqrt(l*w*mult))}
+ nfactor = {1.77182271384+0*(0.02/sqrt(l*w*mult))} wnfactor = 1.93716081040021e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.080000000000001
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.08353125
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0029407877
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 333712830.0
+ pscbe2 = 1.5000958e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 5.0667189e-5
+ alpha1 = 0.0
+ beta0 = 38.266046
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -1.27942399694e-08 wagidl = 1.41921864756822e-13
+ bgidl = 1704700000.0
+ cgidl = -55.9693999999995 wcgidl = 0.0053218703582424
+ egidl = 0.69350825
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.575049627539999 wkt1 = -4.78968332242086e-9
+ kt2 = -0.019032
+ at = 382625.917599999 wat = 0.33350387578319
+ ute = -1.0091712694 wute = -2.65561330876295e-6
+ ua1 = 2.431339464672e-09 wua1 = -1.21420955762801e-14
+ ub1 = -1.8404488054e-18 wub1 = -9.18377428154029e-24
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.34 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.985504201233779+0*(0.0/sqrt(l*w*mult))} lvth0 = 3.17592536828709e-08 wvth0 = 1.02813008558879e-07 pvth0 = 1.28141086030257e-13
+ k1 = 0.604073147499999 lk1 = -6.9793741303501e-8
+ k2 = 0.0192245909377102 lk2 = 8.07156081080825e-09 wk2 = -8.99804271790598e-09 pk2 = 7.89427571287536e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 357633.70352273 lvsat = -1.24130236176009 wvsat = -0.427867466968454 pvsat = 3.36928515538979e-6
+ ua = 2.45225519173184e-09 lua = 1.9985800590439e-15 wua = 1.77443657043906e-18 pua = -4.62823411465753e-23
+ ub = 2.73435708367877e-19 lub = -1.38754965301694e-24 wub = -4.80640047028531e-25 pub = -4.46396454924937e-30
+ uc = -5.147278145e-11 luc = 9.056405360617e-17
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.021419351377321 lu0 = 6.52429670373986e-09 wu0 = -7.61453193117754e-09 pu0 = -1.18263262080749e-14
+ a0 = 0.916336476834248 la0 = -1.85597825970222e-07 wa0 = -1.8081067021916e-08 pa0 = 2.17662586671033e-13
+ keta = -0.00498304443499999 lketa = -2.3173810432149e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.098447303326208 lags = 3.68741832298923e-07 wags = 1.052216220675e-07 pags = -1.19357941474609e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0947625464815+0*(0.009/sqrt(l*w*mult))} lvoff = 1.22677565110199e-8
+ nfactor = {1.89415844162902+0*(0.02/sqrt(l*w*mult))} lnfactor = -9.63344922047457e-07 wnfactor = -6.35384532663913e-07 pnfactor = 6.52883569267299e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.080000000000001
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.641832441643 lpclm = 5.71194892621197e-06 wpclm = -4.2351647362715e-22 ppclm = -6.46234853557053e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 0.004539823205605 lpdiblc2 = -1.25917649924371e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 560098762.7795 lpscbe1 = -1782.69866626545
+ pscbe2 = -1.50486592213e-08 lpscbe2 = 2.36628715770849e-13
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 7.7909598465e-05 lalpha0 = -2.14523077573089e-10
+ alpha1 = 0.0
+ beta0 = 39.13253926505 lbeta0 = -6.82328786496275e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -3.3912576552393e-08 lagidl = 1.66298453256437e-13 wagidl = 2.84821007008082e-13 pagidl = -1.12527358557177e-18
+ bgidl = 1298513669.77135 lbgidl = 3198.55487601853 wbgidl = 1280.1657144237 pbgidl = -0.0100807929348008
+ cgidl = -74.4024181654004 lcgidl = 0.00014515264484526 wcgidl = 0.00707458046389631 pcgidl = -1.38018909979823e-8
+ egidl = 1.2047468705955 legidl = -4.02579964174133e-6
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.608224541233621 lkt1 = 2.61239175371789e-07 wkt1 = 1.62405114011039e-07 pkt1 = -1.31659215108204e-12
+ kt2 = -0.019032
+ at = 710391.088546143 lat = -2.5810196151325 wat = -0.278054483630759 pat = 4.81577745704107e-6
+ ute = -0.47938875450431 lute = -4.17182539179761e-06 wute = -5.2279731402962e-06 pute = 2.02563047293917e-11
+ ua1 = 4.76505314672653e-09 lua1 = -1.83770617607066e-14 wua1 = -2.39035364562438e-14 pua1 = 9.26166423533623e-20
+ ub1 = -4.97533732646125e-19 lub1 = -1.05749190319076e-23 wub1 = -1.49075756167689e-23 pub1 = 4.50726459943912e-29
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.35 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.96115400576174+0*(0.0/sqrt(l*w*mult))} lvth0 = -6.25880136930945e-08 wvth0 = 1.2670682189411e-07 pvth0 = 3.55621168815813e-14
+ k1 = 0.602294036 lk1 = -6.29003958855998e-8
+ k2 = 0.0189935638070392 lk2 = 8.96669853130575e-09 wk2 = 2.96925163768857e-08 pk2 = -7.09676831399267e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -13112.0360914599 lvsat = 0.195189080949051 wvsat = 0.689461964377556 pvsat = -9.59919459303457e-7
+ ua = 3.31666217136051e-09 lua = -1.35065122422537e-15 wua = -2.37606150626435e-17 pua = 5.26557699109291e-23
+ ub = -8.09591033992927e-19 lub = 2.80874576293423e-24 wub = -3.02412203518143e-24 pub = 5.39101076204789e-30
+ uc = -5.44361927e-11 luc = 1.0204608683542e-16
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0226646399527201 lu0 = 1.69930158949885e-09 wu0 = -1.34136316118242e-08 pu0 = 1.06428654145589e-14
+ a0 = 0.818031877417202 la0 = 1.95293174931069e-07 wa0 = 5.60433925882905e-08 pa0 = -6.95400445346858e-14
+ keta = -0.0051939812 lketa = -2.235651484248e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.176526920902361 lags = 6.62145460383608e-08 wags = -2.71794047861343e-07 pags = 2.67205499960204e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0645862731911+0*(0.009/sqrt(l*w*mult))} lvoff = -1.04653231979964e-7
+ nfactor = {1.64013020524995+0*(0.02/sqrt(l*w*mult))} lnfactor = 2.09128826269128e-08 wnfactor = 4.16527313392716e-06 pnfactor = -1.20717925023008e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.0202002600000011 leta0 = 2.31700072604e-7
+ etab = -0.1214502716 letab = 1.9934922234136e-7
+ dsub = 0.810118505 ldsub = -9.69109159472999e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.044838468325 lpclm = -8.23226181550044e-7
+ pdiblc1 = 0.57808555402 lpdiblc1 = -7.28756287605892e-7
+ pdiblc2 = -0.0010893622944 lpdiblc2 = 9.21907714588224e-9
+ pdiblcb = 0.16246 lpdiblcb = -7.26332516e-07 wpdiblcb = -2.11758236813575e-22 ppdiblcb = 2.01948391736579e-28
+ drout = 0.147588000000001 ldrout = 1.5979315352e-6
+ pscbe1 = -151521249.434 lpscbe1 = 974.544233056977
+ pscbe2 = 7.55293005675e-08 lpscbe2 = -1.14324647226836e-13
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 4.36726325897e-05 lalpha0 = -8.18685295926516e-11
+ alpha1 = -9.37299999999999e-11 lalpha1 = 3.63166258e-16
+ beta0 = 69.5879243857 lbeta0 = -0.000124825723053433
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.66790829307034e-08 lagidl = -2.97239905767686e-14 wagidl = -5.27970752101699e-14 pagidl = 1.8286143579107e-19
+ bgidl = 2971288240.4573 lbgidl = -3282.77747556126 wbgidl = -2560.33142884738 pbgidl = 0.0047995972965173
+ cgidl = -510.735397289199 lcgidl = 0.00183576840575833 wcgidl = 0.00680463923371518 pcgidl = -1.27559767075225e-8
+ egidl = -1.553543708466 legidl = 6.66147303589036e-06 wegidl = 8.470329472543e-22 pegidl = 4.8467614016779e-27
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.54173832 lkt1 = 3.63166258000002e-09 wkt1 = -1.77395678608078e-7
+ kt2 = -0.019032
+ at = -164261.409914206 lat = 0.80790895540197 wat = 2.63406943735569 pat = -6.46753788721304e-6
+ ute = -1.82003516969092 lute = 1.02264320848444e-06 wute = 8.28039388405575e-07 pute = -3.20832141431626e-12
+ ua1 = -4.749579392e-10 lua1 = 1.92588519282432e-15 wua1 = -6.90253292068385e-31 pua1 = 2.44502824971036e-36
+ ub1 = -2.64869845781944e-18 lub1 = -2.24001618775111e-24 wub1 = -7.53796316660695e-24 pub1 = 1.65183455949937e-29
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.36 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.0970119945346+0*(0.0/sqrt(l*w*mult))} lvth0 = 1.92091372060505e-07 wvth0 = 5.74573159925932e-07 pvth0 = -8.04008120392862e-13
+ k1 = 0.55942551 lk1 = 1.74609429539999e-8
+ k2 = 0.00913940723257972 lk2 = 2.74393004457876e-08 wk2 = 5.61949056165057e-08 pk2 = -1.20649062008518e-13
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 128725.538692 lvsat = -0.0706996367400233 wvsat = 0.332545939118707 pvsat = -2.90844678353221e-7
+ ua = 3.42594614659591e-09 lua = -1.55551496420166e-15 wua = -1.10593482794107e-17 pua = 2.88459751990691e-23
+ ub = 2.24322915843054e-18 lub = -2.91407096978279e-24 wub = -1.09843072818996e-23 pub = 2.03131740255457e-29
+ uc = 5.12043316e-13 luc = -9.59876400173601e-19
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0319932082351523 lu0 = -1.57880325127487e-08 wu0 = -3.71804868335447e-08 pu0 = 5.5196212213196e-14
+ a0 = 1.05037937213657 la0 = -2.40265438669851e-07 wa0 = -2.68017070451665e-07 pa0 = 5.37943699480008e-13
+ keta = 0.0419609792 lketa = -1.1075320360832e-07 pketa = -1.0097419586829e-28
+ a1 = 0.0
+ a2 = 0.5
+ ags = -0.170448996413385 lags = 7.16655600638457e-07 wags = -7.41666250640175e-07 pags = 1.1480279312894e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.2251322265544+0*(0.009/sqrt(l*w*mult))} lvoff = 1.96306212194878e-07 wvoff = 4.74558101823854e-07 pvoff = -8.89606617678997e-13
+ nfactor = {1.0623624380501+0*(0.02/sqrt(l*w*mult))} lnfactor = 1.10399633901974e-06 wnfactor = -9.14963412840077e-07 pnfactor = -2.54838107173092e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.4373e-05 lcit = -8.1976258e-12
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.270598149321284 leta0 = -2.37695810717677e-07 weta0 = -7.51502868337964e-09 peta0 = 1.40876727698624e-14
+ etab = -0.0283214568 letab = 2.476994611728e-8
+ dsub = -0.466714193220436 ldsub = 1.42444141661103e-06 wdsub = 3.80381893693904e-06 pdsub = -7.13063897918592e-12
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.0831858186719989 lpclm = 9.7948787548947e-7
+ pdiblc1 = 0.00549710251999991 lpdiblc1 = 3.44618023576008e-7
+ pdiblc2 = 0.00585964945018 lpdiblc2 = -3.80754027050743e-9
+ pdiblcb = -0.39992 lpdiblcb = 3.27905032e-07 ppdiblcb = 8.07793566946316e-28
+ drout = 1.515411042014 ldrout = -9.66189539359445e-7
+ pscbe1 = 428577028.488 lpscbe1 = -112.907998735605
+ pscbe2 = 1.45331535696e-08 lpscbe2 = 1.87299354278326e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -5.93092031506e-05 lalpha0 = 1.11181219686115e-10 walpha0 = -7.1131193393326e-26 palpha0 = -9.74486697622638e-32
+ alpha1 = 1.8746e-10 lalpha1 = -1.63952516e-16
+ beta0 = -38.239948205 lbeta0 = 7.7308406905093e-05 wbeta0 = -4.06575814682064e-20
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -3.71324370668416e-09 lagidl = 8.50346493767805e-15 wagidl = 6.94994034423295e-14 pagidl = -4.63955430909058e-20
+ bgidl = 534379280.870919 lbgidl = 1285.45206007937 wbgidl = 1940.92975898794 pbgidl = -0.0036384669261988
+ cgidl = 556.49103 lcgidl = -0.000164854254838
+ egidl = 3.067904826664 legidl = -2.00189438806434e-6
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.460912992092 lkt1 = -1.47883497116337e-07 wkt1 = -3.32545939118707e-07 pkt1 = 2.90844678353222e-13
+ kt2 = -0.019032
+ at = 473746.5163768 lat = -0.388100703223149 wat = -1.52971131994605 pat = 1.33788552042482e-6
+ ute = -1.11157904061816 lute = -3.05428651075357e-07 wute = -1.65607877681116e-06 pute = 1.44840649819905e-12
+ ua1 = 5.524e-10
+ ub1 = -4.06466517677944e-18 lub1 = 4.14355023611299e-25 wub1 = 2.38767984287232e-24 pub1 = -2.08826479057612e-30
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.81e-6
+ sbref = 2.81e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.37 pmos
* DC IV MOS Parameters
+ lmin = 8.0e-07 lmax = 1e-06 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.676228052033682+0*(0.0/sqrt(l*w*mult))} lvth0 = -1.75926264050794e-07 wvth0 = -1.99186088675415e-06 pvth0 = 1.44059509683353e-12
+ k1 = 0.589711379999999 lk1 = -9.02707894799971e-9
+ k2 = 0.0582594263814829 lk2 = -1.55210683018431e-08 wk2 = -3.20466774659412e-07 pk2 = 2.087792435608e-13
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 8829.08188871259 lvsat = 0.034161804380132 wvsat = 0.0238205373892524 pvsat = -2.08334420006402e-8
+ ua = -7.19970537316832e-10 lua = 2.07050376754843e-15 wua = 1.49561386239831e-16 pua = -1.11632919211451e-22
+ ub = -3.92188615630164e-18 lub = 2.47793888448196e-24 wub = 5.40460802205743e-23 pub = -3.65624028841179e-29
+ uc = 5.75692682e-12 luc = -5.547051512772e-18 puc = -5.87747175411144e-39
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = -0.00222669788070629 lu0 = 1.41406973761813e-08 wu0 = 1.22126784252487e-07 pu0 = -8.41339270786473e-14
+ a0 = 0.546822571003945 la0 = 2.00145339600738e-07 wa0 = 1.51767984831494e-06 pa0 = -1.02382682567326e-12
+ keta = -0.150384786 lketa = 5.74724026356e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.405566781876555 lags = 2.12872200946075e-07 wags = 2.49683314239752e-06 pags = -1.68436363786137e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {0.242654183714998+0*(0.009/sqrt(l*w*mult))} lvoff = -2.12819782226738e-07 wvoff = -2.37279050911927e-06 pvoff = 1.60068447745186e-12
+ nfactor = {3.53478033742152+0*(0.02/sqrt(l*w*mult))} lnfactor = -1.0583803557705e-06 wnfactor = -1.42329385205548e-05 pnfactor = 9.09951995747636e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -1.1865e-05 lcit = 1.4750129e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.00021886458217845 leta0 = -1.22208828485498e-09 weta0 = -1.59584849129217e-09 peta0 = 8.91075777386342e-15
+ etab = -0.0019949792217191 letab = 1.74480882731552e-09 wetab = 1.90965197382064e-08 petab = -1.67018161630353e-14
+ dsub = 4.15432788975418 ldsub = -2.61712198915857e-06 wdsub = -1.90193047075192e-05 pdsub = 1.28304649602572e-11
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.98195455905 lpclm = -6.8117526484513e-7
+ pdiblc1 = 0.20581194057 lpdiblc1 = 1.69422666217479e-7
+ pdiblc2 = -0.0319025077049 lpdiblc2 = 2.92192423773255e-08 wpdiblc2 = -2.64697796016969e-23 ppdiblc2 = -3.78653234506086e-29
+ pdiblcb = -0.025
+ drout = 0.33949907438 ldrout = 6.22630675332523e-8
+ pscbe1 = -39572648.1000004 lpscbe1 = 296.53570840826
+ pscbe2 = 1.8099436842e-08 lpscbe2 = -3.10034141461322e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.00023839585627 lalpha0 = -1.49191625283142e-10
+ alpha1 = 0.0
+ beta0 = 66.364220735 lbeta0 = -1.4178399249831e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 3.34009768491444e-08 lagidl = -2.39566323604496e-14 wagidl = -2.47937740762248e-13 pagidl = 2.31234983230417e-19
+ bgidl = 2668077995.6454 lbgidl = -580.680835862386 wbgidl = -9704.6487949397 pbgidl = 0.00654675607706631
+ cgidl = -144.696 lcgidl = 0.000448403921599999
+ egidl = 1.78393816687 legidl = -8.78937147408502e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.558965652137999 lkt1 = -6.21266406401052e-08 wkt1 = -1.79506687183516e-07 pkt1 = 1.56996548610701e-13
+ kt2 = -0.019032
+ at = 46865.0 lat = -0.014750129
+ ute = -1.396713 lute = -5.60504902000005e-8
+ ua1 = 5.524e-10
+ ub1 = -3.5909e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.41e-6
+ sbref = 2.41e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.38 pmos
* DC IV MOS Parameters
+ lmin = 6e-07 lmax = 8.0e-07 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.935543057763581+0*(0.0/sqrt(l*w*mult))} lvth0 = -9.92361185403865e-10 wvth0 = 4.8442871314592e-07 pvth0 = -2.29909867259052e-13
+ k1 = 0.593154569999998 lk1 = -1.13498549220005e-8
+ k2 = 0.020870327675526 lk2 = 9.70161768519534e-09 wk2 = -3.70382131221987e-08 pk2 = 1.75783359477956e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 63090.3015112873 lvsat = -0.00244281437725696 wvsat = -0.0238205373892524 pvsat = 1.13052270449391e-8
+ ua = -1.72654669752753e-09 lua = 2.74954004522657e-15 wua = -5.36940402703154e-17 pua = 2.54831915122987e-23
+ ub = 2.5023217714044e-18 lub = -1.85583178354853e-24 wub = -5.14585836592746e-25 pub = 2.44222438046917e-31
+ uc = 2.42542760000001e-12 luc = -3.29962213896e-18
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.00877686002928396 lu0 = 6.71769721010183e-09 wu0 = -8.73599210959773e-09 pu0 = 4.14610185521517e-15
+ a0 = 0.932568689999998 la0 = -6.00789922740004e-8
+ keta = 0.0100696950000002 lketa = -5.0770190247e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = -0.533912240000001 lags = 8.46644749104e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {0.00559779755700007+0*(0.009/sqrt(l*w*mult))} lvoff = -5.29015441245522e-8
+ nfactor = {2.1244191892703+0*(0.02/sqrt(l*w*mult))} lnfactor = -1.06950725227682e-07 wnfactor = -2.51010184244951e-06 pnfactor = 1.19129433442654e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -0.0616384141885894 leta0 = 4.0506831973905e-08 weta0 = 3.91709919081887e-08 peta0 = -1.85905527596263e-14
+ etab = 0.0019949792217191 letab = -9.46817138627884e-10 wetab = -1.90965197382064e-08 petab = 9.06320826775275e-15
+ dsub = 0.195107531568001 ldsub = 5.37680644738264e-08 wdsub = 2.10022824001857e-10 pdsub = -9.9676832273097e-17
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.272763882949999 lpclm = 4.7184476525193e-7
+ pdiblc1 = 0.195445235049998 lpdiblc1 = 1.7641604576127e-7
+ pdiblc2 = 0.0256746597612 lpdiblc2 = -9.62231479530552e-9
+ pdiblcb = -0.025
+ drout = -0.658708114820001 ldrout = 7.35653637367572e-7
+ pscbe1 = 430031833.719999 lpscbe1 = -20.2594750275121
+ pscbe2 = 1.0746893781e-08 lpscbe2 = 1.85968413433739e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -0.000112188837415 lalpha0 = 8.73128090767591e-11 walpha0 = -2.06795153138257e-25 palpha0 = 9.86076131526265e-32
+ alpha1 = 0.0
+ beta0 = 27.750617018 lbeta0 = 1.18703378176572e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -2.2596237190084e-08 lagidl = 1.38190882304139e-14 wagidl = 3.19880916561026e-13 pagidl = -1.51815482999863e-19
+ bgidl = 2044837300 lbgidl = -160.242662579998
+ cgidl = 1208.17 lcgidl = -0.000464239482
+ egidl = -0.197226229600001 legidl = 4.5755635445016e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.728371307861998 lkt1 = 5.21544147113049e-08 wkt1 = 1.79506687183516e-07 pkt1 = -8.51938737372977e-14
+ kt2 = -0.019032
+ at = 41610.9999999999 lat = -0.0112057806
+ ute = -1.6043825 lute = 8.40433545000009e-8
+ ua1 = 5.53349199999999e-10 lua1 = -6.40330320000131e-19
+ ub1 = -4.2831041e-18 lub1 = 4.6696088586e-25
+ uc1 = -2.69861592e-10 luc1 = 1.083823099632e-16 puc1 = 3.76158192263132e-37
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.02e-6
+ sbref = 2.01e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.39 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 6e-07 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.06103555822525+0*(0.0/sqrt(l*w*mult))} lvth0 = 5.85663795337052e-08 wvth0 = 1.08111444060995e-06 pvth0 = -5.13096913513489e-13
+ k1 = 0.351195792613638 lk1 = 1.03483780825567e-07 wk1 = 7.75499755480873e-07 pk1 = -3.68052183951224e-13
+ k2 = 0.0192423241922279 lk2 = 1.04742681383686e-08 wk2 = 9.69540825404106e-08 pk2 = -4.60144075736789e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 97450.2129484891 lvsat = -0.0187500283453529 wvsat = -0.403273163334294 pvsat = 1.91393443318456e-7
+ ua = 1.75664231131689e-08 lua = -6.40690342692994e-15 wua = -4.4732243326281e-14 pua = 2.12299226826529e-20
+ ub = -6.43891241843284e-18 lub = 2.38767796294823e-24 wub = -5.26768342904616e-24 pub = 2.5000425554253e-30
+ uc = -4.48034609955098e-11 luc = 1.91152083884689e-17 wuc = 3.03435045713518e-16 puc = -1.44010272695635e-22
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0656613693046714 lu0 = -2.0279690891997e-08 wu0 = -1.79514570647474e-07 pu0 = 8.51976152292912e-14
+ a0 = -1.28760245098549 la0 = 9.93614231237713e-07 wa0 = 1.06862138542313e-05 pa0 = -5.07167709521815e-12
+ keta = -0.0417133953527917 lketa = -2.6193935565565e-08 wketa = -6.79542459258559e-07 pketa = 3.22510851164112e-13
+ a1 = 0.0
+ a2 = 0.5
+ ags = 1.25
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.418673339105244+0*(0.009/sqrt(l*w*mult))} lvoff = 1.48457537335349e-07 wvoff = 2.08787526713188e-06 pvoff = -9.90905601780789e-13
+ nfactor = {-5.84315913056827+0*(0.02/sqrt(l*w*mult))} lnfactor = 3.6744619453677e-06 wnfactor = 4.98911487934814e-05 pnfactor = -2.36783392173863e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 2.873e-05 lcit = -8.88925800000001e-12 wcit = 1.03397576569128e-25
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -0.562367586009025 leta0 = 2.78152896919884e-07 weta0 = 2.64002178969529e-06 peta0 = -1.25295434138938e-12
+ etab = -0.0457887566537599 letab = 2.17313439078744e-08 wetab = 4.23880059150457e-07 petab = -2.01173476072807e-13
+ dsub = 0.518144002163548 ldsub = -9.95450444708201e-08 wdsub = -7.18952067655127e-07 pdsub = 3.41214651309124e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.433002908249321 lpclm = 8.06801684355126e-07 wpclm = 1.01300137339743e-05 ppclm = -4.80770451814418e-12
+ pdiblc1 = 2.52162806827304 lpdiblc1 = -9.27590326886382e-07 wpdiblc1 = -6.55631814869689e-06 ppdiblc1 = 3.11162859337155e-12
+ pdiblc2 = 0.0375524862945939 lpdiblc2 = -1.52595312680543e-08 wpdiblc2 = -2.10544847701512e-07 ppdiblc2 = 9.99245847191375e-14
+ pdiblcb = -0.025
+ drout = -0.809838006837193 ldrout = 8.07379884118931e-07 wdrout = 1.17580575175587e-05 pdrout = -5.58037409783335e-12
+ pscbe1 = 54569310.9023476 lpscbe1 = 157.935038301746 wpscbe1 = 2994.15006492625 ppscbe1 = -0.001421023620814
+ pscbe2 = 1.50747496741437e-08 lpscbe2 = -1.94316272548606e-16 wpscbe2 = 1.82724222591753e-15 ppscbe2 = -8.67209160420406e-22
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -0.000523993688909691 lalpha0 = 2.82755391596139e-10 walpha0 = 3.52556177076268e-09 palpha0 = -1.67323161640397e-15
+ alpha1 = 0.0
+ beta0 = 6.38109055790721 lbeta0 = 2.20123150756172e-05 wbeta0 = 0.000275808913550145 pbeta0 = -1.30898910370899e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 6.27623796007204e-09 lagidl = 1.16211524149804e-16 wagidl = -9.52927720102458e-14 pagidl = 4.52259495960626e-20
+ bgidl = 3350871044.25681 lbgidl = -780.08627760428 wbgidl = -7615.44747027487 pbgidl = 0.00361429136939245
+ cgidl = 2573.11156720801 lcgidl = -0.00111204074979692 wcgidl = -0.0150182471926887 pcgidl = 7.12766011765004e-9
+ egidl = 1.23295061677587 legidl = -2.21205576839826e-07 wegidl = -6.02040329453731e-07 pegidl = 2.85728340358746e-13
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.485879241839999 lkt1 = -6.29323198227365e-08 wkt1 = -1.32904842413174e-06 pkt1 = 6.30766382092924e-13
+ kt2 = -0.019032
+ at = 18000.0
+ ute = -1.6329554 lute = 9.76040528399988e-8
+ ua1 = 5.52e-10
+ ub1 = -1.4495264024472e-17 lub1 = 5.31365198601443e-24 wub1 = 4.87760771656349e-23 pub1 = -2.31491262228103e-29
+ uc1 = -4.1496e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 1.81e-6
+ sbref = 1.81e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.40 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.982438509334+0*(0.0/sqrt(l*w*mult))} wvth0 = 1.23961389355456e-7
+ k1 = 0.59521
+ k2 = 0.02024257534638 wk2 = 1.06236205213546e-9
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200000.0
+ ua = 2.70553474874766e-09 wua = -1.47584754910791e-18
+ ub = -1.74654515799999e-20 wub = -4.69479920508922e-25
+ uc = -3.9972e-11
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0214495801802 wu0 = -5.09311794985126e-9
+ a0 = 0.892355895310459 wa0 = 1.16334351390839e-8
+ keta = -0.0079259
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.150195232522 wags = -7.11535157710457e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.093204657+0*(0.009/sqrt(l*w*mult))}
+ nfactor = {1.80413481106+0*(0.02/sqrt(l*w*mult))} wnfactor = 3.08697027190568e-8
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.080000000000001
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.08353125
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0029407877
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 333712830.0
+ pscbe2 = 1.5000958e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 5.0667189e-5
+ alpha1 = 0.0
+ beta0 = 38.266046
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.6264259718e-08 wagidl = -4.52704573373753e-15
+ bgidl = 1596787242.0 wbgidl = 543.858286117365
+ cgidl = 1000.0
+ egidl = 0.69350825
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.576
+ kt2 = -0.019032
+ at = 448800.0
+ ute = -1.5361
+ ua1 = 2.2096e-11
+ ub1 = -3.6627e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.41 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.982438509334+0*(0.0/sqrt(l*w*mult))} wvth0 = 1.23961389355454e-7
+ k1 = 0.59521
+ k2 = 0.02024257534638 wk2 = 1.06236205213549e-9
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200000.0
+ ua = 2.70553474874766e-09 wua = -1.47584754910791e-18
+ ub = -1.746545158e-20 wub = -4.69479920508922e-25
+ uc = -3.9972e-11
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0214495801802 wu0 = -5.09311794985124e-9
+ a0 = 0.892355895310459 wa0 = 1.16334351390856e-8
+ keta = -0.0079259
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.150195232522 wags = -7.11535157710455e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.093204657+0*(0.009/sqrt(l*w*mult))}
+ nfactor = {1.80413481106+0*(0.02/sqrt(l*w*mult))} wnfactor = 3.08697027190568e-8
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.080000000000001
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.08353125
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0029407877
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 333712830.0
+ pscbe2 = 1.5000958e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 5.0667189e-5
+ alpha1 = 0.0
+ beta0 = 38.266046
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.6264259718e-08 wagidl = -4.52704573373753e-15
+ bgidl = 1596787242.0 wbgidl = 543.858286117367
+ cgidl = 1000.0
+ egidl = 0.69350825
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.576
+ kt2 = -0.019032
+ at = 448800.0
+ ute = -1.5361
+ ua1 = 2.2096e-11
+ ub1 = -3.6627e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.42 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.992159134544159+0*(0.0/sqrt(l*w*mult))} lvth0 = 7.65460352799159e-08 wvth0 = 1.363525148368e-07 pvth0 = -9.75751567153908e-14
+ k1 = 0.6040731475 lk1 = -6.9793741303501e-8
+ k2 = 0.0161389483980739 lk2 = 3.23144207671306e-08 wk2 = 6.55296621078232e-09 pk2 = -4.32363115076806e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 272735.9285 lvsat = -0.5727663425661
+ ua = 2.45253548351987e-09 lua = 1.99226801396278e-15 wua = 3.61823138298062e-19 pua = -1.44709215950102e-23
+ ub = 3.32702434415952e-19 lub = -2.75743203506372e-24 wub = -7.79332255898715e-25 pub = 2.43996320026047e-30
+ uc = -5.147278145e-11 luc = 9.056405360617e-17
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0211203070405256 lu0 = 2.59289426568008e-09 wu0 = -6.10740947877327e-09 pu0 = 7.9871400736495e-15
+ a0 = 0.909308152606532 la0 = -1.33492245303655e-07 wa0 = 1.73402533076289e-08 pa0 = -4.49389103500055e-14
+ keta = -0.004983044435 lketa = -2.3173810432149e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.138085641377428 lags = 9.53581864270445e-08 wags = -9.45475154896873e-08 pags = 1.84218390184416e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0947625464815+0*(0.009/sqrt(l*w*mult))} lvoff = 1.22677565110199e-8
+ nfactor = {1.71068135050411+0*(0.02/sqrt(l*w*mult))} lnfactor = 7.35908620493426e-07 wnfactor = 2.89302577279079e-07 pnfactor = -2.03505551401034e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.080000000000001
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.641832441643001 lpclm = 5.71194892621197e-06 wpclm = 2.11758236813575e-22 ppclm = 3.23117426778526e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 0.004539823205605 lpdiblc2 = -1.25917649924371e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 560098762.7795 lpscbe1 = -1782.69866626545
+ pscbe2 = -1.50486592213e-08 lpscbe2 = 2.36628715770849e-13
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 7.7909598465e-05 lalpha0 = -2.14523077573089e-10
+ alpha1 = 0.0
+ beta0 = 39.13253926505 lbeta0 = -6.82328786496275e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 2.65844372871815e-08 lagidl = -8.12672702862767e-14 wagidl = -2.00716013525502e-14 pagidl = 1.22407157675902e-19
+ bgidl = 1340082633.9633 lbgidl = 2021.4461064458 wbgidl = 1070.66661496496 pbgidl = -0.00414840486634321
+ cgidl = 1329.341 lcgidl = -0.0025934286386 wcgidl = -1.73472347597681e-18
+ egidl = 1.2047468705955 legidl = -4.02579964174133e-06 pegidl = 6.46234853557053e-27
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.576
+ kt2 = -0.019032
+ at = 646326.929845892 lat = -1.55544556176446 wat = 0.0448158071301332 pat = -3.52906554826944e-7
+ ute = -1.516727 lute = -1.525546258e-7
+ ua1 = 2.2096e-11
+ ub1 = -3.2744191136829e-18 lub1 = -3.05755666739264e-24 wub1 = -9.12639780961318e-25 pub1 = 7.18667321915798e-30
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.43 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.953644791945492+0*(0.0/sqrt(l*w*mult))} lvth0 = -7.26816365528779e-08 wvth0 = 8.88619161398464e-08 pvth0 = 8.64319169958231e-14
+ k1 = 0.602294036 lk1 = -6.29003958855998e-8
+ k2 = 0.0285006729392287 lk2 = -1.55823171400273e-08 wk2 = -1.82213741990859e-08 pk2 = 5.27543478443948e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 137937.513954 lvsat = -0.0504764055661682 wvsat = -0.0717969537433532 pvsat = 2.78184476973997e-7
+ ua = 3.31344302741963e-09 lua = -1.34340435563123e-15 wua = -7.53678630594257e-18 pua = 1.61330305576124e-23
+ ub = -1.42713869215565e-18 lub = 4.0612483939506e-24 wub = 8.81921822364053e-26 pub = -9.21346987737879e-31
+ uc = -5.44361927e-11 luc = 1.0204608683542e-16
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0202440735996622 lu0 = 5.98794835564961e-09 wu0 = -1.21447098794838e-09 pu0 = -1.09710394029005e-14
+ a0 = 0.828819013815985 la0 = 1.78370971854204e-07 wa0 = 1.67842571424984e-09 pa0 = 1.57444068432969e-14
+ keta = -0.00519398120000001 lketa = -2.235651484248e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.127255035752035 lags = 1.37322450983194e-07 wags = -2.34737981682698e-08 pags = -9.11638349491486e-14
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0645862731911001+0*(0.009/sqrt(l*w*mult))} lvoff = -1.04653231979964e-7
+ nfactor = {2.77484801695985+0*(0.02/sqrt(l*w*mult))} lnfactor = -3.38731154535601e-06 wnfactor = -1.55347315465716e-06 pnfactor = 5.10496333694982e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.020200260000001 leta0 = 2.31700072604e-7
+ etab = -0.1214502716 letab = 1.9934922234136e-7
+ dsub = 0.810118505 ldsub = -9.69109159473e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.04483730015268 lpclm = -8.23221655349557e-07 wpclm = 5.88735020648067e-12 ppclm = -2.28111271110524e-17
+ pdiblc1 = 0.57808555402 lpdiblc1 = -7.28756287605892e-7
+ pdiblc2 = -0.0010893622944 lpdiblc2 = 9.21907714588224e-9
+ pdiblcb = 0.16246 lpdiblcb = -7.26332516e-07 wpdiblcb = -5.29395592033938e-23
+ drout = 0.147588000000001 ldrout = 1.5979315352e-6
+ pscbe1 = -151521249.434 lpscbe1 = 974.544233056976
+ pscbe2 = 7.55293005675e-08 lpscbe2 = -1.14324647226836e-13
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 4.36726325897e-05 lalpha0 = -8.18685295926516e-11
+ alpha1 = -9.37299999999999e-11 lalpha1 = 3.63166258e-16
+ beta0 = 69.5879243857 lbeta0 = -0.000124825723053433
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.22163573986367e-09 lagidl = 1.70034405889611e-14 wagidl = 2.51053053124351e-14 pagidl = -5.26352848882499e-20
+ bgidl = 2463265410.0 lbgidl = -2330.437877586 wbgidl = 3.63797880709171e-12
+ cgidl = 839.446085 lcgidl = -0.000695281800941
+ egidl = -1.553543708466 legidl = 6.66147303589036e-06 wegidl = 4.2351647362715e-22 pegidl = -1.61558713389263e-27
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.5769373 lkt1 = 3.63166258000002e-9
+ kt2 = -0.019032
+ at = 471525.844772338 lat = -0.878161277538469 wat = -0.57016862566453 pat = 2.02991212847926e-6
+ ute = -1.65573499 lute = 3.86045732254e-7
+ ua1 = -4.749579392e-10 lua1 = 1.92588519282432e-15 wua1 = -4.93038065763132e-32 pua1 = 1.50463276905253e-36
+ ub1 = -5.26288026255206e-18 lub1 = 4.64693490001581e-24 wub1 = 5.63697983615726e-24 pub1 = -1.81904829493297e-29
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.44 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.976938432589611+0*(0.0/sqrt(l*w*mult))} lvth0 = -2.90153778014112e-08 wvth0 = -3.05730972701589e-08 pvth0 = 3.10324793134222e-13
+ k1 = 0.55942551 lk1 = 1.74609429539999e-8
+ k2 = 0.0229722191732166 lk2 = -5.21867771026116e-09 wk2 = -1.35196446706685e-08 pk2 = 4.39404856704236e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 166217.538692 lvsat = -0.103490139940023 wvsat = 0.143593907486707 pvsat = -1.25587231487874e-7
+ ua = 3.42088585113187e-09 lua = -1.5448166729622e-15 wua = 1.44435085591058e-17 pua = -2.50712301963887e-23
+ ub = -7.54259685597031e-19 lub = 2.79986940825582e-24 wub = 4.12242500427521e-24 pub = -8.48391983593182e-30
+ uc = 5.12043316e-13 luc = -9.59876400173601e-19
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0240036176606338 lu0 = -1.05969294104781e-09 wu0 = 3.08541978555182e-09 pu0 = -1.90316146469039e-14
+ a0 = 0.985633276640952 la0 = -1.15593045237482e-07 wa0 = 5.82900426427506e-08 pa0 = -9.03797302508683e-14
+ keta = 0.0419609792 lketa = -1.1075320360832e-07 pketa = -2.52435489670724e-29
+ a1 = 0.0
+ a2 = 0.5
+ ags = -0.385603260112601 lags = 1.09872661241104e-06 wags = 3.42667346934079e-07 pags = -7.77532025558011e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0903106772300004+0*(0.009/sqrt(l*w*mult))} lvoff = -5.64302641686413e-08 wvoff = -2.04915003175055e-07 pvoff = 3.8413366495196e-13
+ nfactor = {0.768973129903674+0*(0.02/sqrt(l*w*mult))} lnfactor = 3.72901517919502e-07 wnfactor = 5.63658848799056e-07 pnfactor = 1.13618768327079e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.4373e-05 lcit = -8.1976258e-12
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.280071646278664 leta0 = -2.55454828113981e-07 weta0 = -5.52595207551953e-08 peta0 = 1.03589497607689e-13
+ etab = -0.0283214568 letab = 2.476994611728e-8
+ dsub = 0.288041671348605 ldsub = 9.57607288990563e-09 wdsub = 3.34970744379575e-12 pdsub = -6.27936157431935e-18
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.0831881550166482 lpclm = 9.7948583212244e-07 wpclm = -1.17747004146554e-11 ppclm = 1.02981529827238e-17
+ pdiblc1 = 0.00549710251999969 lpdiblc1 = 3.44618023576008e-7
+ pdiblc2 = 0.00585964945018 lpdiblc2 = -3.80754027050743e-9
+ pdiblcb = -0.39992 lpdiblcb = 3.27905032e-07 wpdiblcb = -4.2351647362715e-22
+ drout = 1.515411042014 ldrout = -9.66189539359445e-07 wdrout = -1.6940658945086e-21
+ pscbe1 = 428577028.488 lpscbe1 = -112.907998735605
+ pscbe2 = 1.45331535696e-08 lpscbe2 = 1.87299354278579e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -5.93092031506001e-05 lalpha0 = 1.11181219686115e-10 walpha0 = -2.82806634521733e-28 palpha0 = 1.26592278024234e-32
+ alpha1 = 1.8746e-10 lalpha1 = -1.63952516e-16
+ beta0 = -38.239948205 lbeta0 = 7.73084069050931e-05 wbeta0 = 2.03287907341032e-20 pbeta0 = -1.93870456067116e-26
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 6.84992395057597e-09 lagidl = 6.45265150915977e-15 wagidl = 1.62631933359405e-14 pagidl = -3.60598617771132e-20
+ bgidl = 919499980.0 lbgidl = 563.504797492001
+ cgidl = 1290.2661705216 lcgidl = -0.00154038913325979 wcgidl = -0.0036980770181002 pcgidl = 6.93241517813063e-9
+ egidl = 3.067904826664 legidl = -2.00189438806434e-6
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.526897 lkt1 = -9.01738838e-8
+ kt2 = -0.019032
+ at = -20476.9289282439 lat = 0.0441471220406421 wat = 0.961074022808528 pat = -8.40555340348339e-7
+ ute = -1.4401794 lute = -1.80347767599999e-8
+ ua1 = 5.524e-10
+ ub1 = -2.07825930016428e-18 lub1 = -1.32295555607632e-24 wub1 = -7.62340054846926e-24 pub1 = 6.66742611969121e-30
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.81e-6
+ sbref = 2.81e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.45 pmos
* DC IV MOS Parameters
+ lmin = 8.0e-07 lmax = 1e-06 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.35280081372142+0*(0.0/sqrt(l*w*mult))} lvth0 = 2.99713860736474e-07 wvth0 = 1.4179278113087e-06 pvth0 = -9.56534101508844e-13
+ k1 = 0.58971138 lk1 = -9.02707894799971e-9
+ k2 = -0.0371904285068295 lk2 = 4.73995739507071e-08 wk2 = 1.60581022207285e-07 pk2 = -1.08327957581034e-13
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 13555.5703 lvsat = 0.03002801761562
+ ua = -6.77953742531332e-10 lua = 2.04002843565564e-15 wua = -6.21946880529614e-17 pua = 4.19565365605256e-23
+ ub = 1.16419015161633e-17 lub = -8.04181317880374e-24 wub = -2.43922346359636e-23 pub = 1.64550014854211e-29
+ uc = 5.75692682e-12 luc = -5.547051512772e-18 wuc = -3.08148791101958e-33 puc = 1.46936793852786e-39
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0382099223247124 lu0 = -1.3484527000251e-08 wu0 = -8.16655325123017e-08 pu0 = 5.50915682327987e-14
+ a0 = 0.887049862563472 la0 = -2.93719912853178e-08 wa0 = -1.969962947776e-07 pa0 = 1.32893700456969e-13
+ keta = -0.150384786 lketa = 5.74724026355999e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 1.37505224558279 lags = -4.41142692870154e-07 wags = -2.38917581964733e-06 pags = 1.61173800793409e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.431453562906998+0*(0.009/sqrt(l*w*mult))} lvoff = 2.41933303644461e-07 wvoff = 1.02457501587528e-06 pvoff = -6.91178305709463e-13
+ nfactor = {-0.90562897333372+0*(0.02/sqrt(l*w*mult))} lnfactor = 1.83750851741093e-06 wnfactor = 8.14581856215223e-06 pnfactor = -5.49516920202789e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -1.1865e-05 lcit = 1.4750129e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -0.0549209570033122 leta0 = 3.75297027164351e-08 weta0 = 2.76297603775977e-07 peta0 = -1.86390363507274e-13
+ etab = 0.00179416616 letab = -1.569177723536e-9
+ dsub = 0.380506894026977 ldsub = -7.12940108645984e-08 wdsub = -1.67485372172847e-11 pdsub = 1.12985632075316e-17
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.98195455905 lpclm = -6.8117526484513e-7
+ pdiblc1 = 0.205811940569999 lpdiblc1 = 1.69422666217478e-7
+ pdiblc2 = -0.0319025077049 lpdiblc2 = 2.92192423773255e-08 ppdiblc2 = -6.31088724176809e-30
+ pdiblcb = -0.025
+ drout = 0.339499074379999 ldrout = 6.22630675332519e-8
+ pscbe1 = -39572648.1000004 lpscbe1 = 296.53570840826
+ pscbe2 = 1.8099436842e-08 lpscbe2 = -3.10034141461322e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.00023839585627 lalpha0 = -1.49191625283142e-10 palpha0 = 1.97215226305253e-31
+ alpha1 = 0.0
+ beta0 = 66.3642207349999 lbeta0 = -1.41783992498309e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 5.86863698166759e-09 lagidl = 7.31088509216701e-15 wagidl = -1.09180364427498e-13 pagidl = 7.36530738427903e-20
+ bgidl = 742474500.0 lbgidl = 718.3312823
+ cgidl = -3813.571702608 lcgidl = 0.00292342747057936 wcgidl = 0.018490385090501 pcgidl = -1.2473613782052e-8
+ egidl = 1.78393816687 legidl = -8.78937147408502e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.594583500000001 lkt1 = -3.09752709000001e-8
+ kt2 = -0.019032
+ at = 46864.9999999999 lat = -0.014750129
+ ute = -1.396713 lute = -5.60504901999988e-8
+ ua1 = 5.524e-10
+ ub1 = -3.5909e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.41e-6
+ sbref = 2.41e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.46 pmos
* DC IV MOS Parameters
+ lmin = 6e-07 lmax = 8.0e-07 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.617208859136104+0*(0.0/sqrt(l*w*mult))} lvth0 = -1.96516471826783e-07 wvth0 = -1.11991070776005e-06 pvth0 = 7.55491763454932e-13
+ k1 = 0.618726200293859 lk1 = -2.86004767182378e-08 wk1 = -1.28875800068475e-07 pk1 = 8.69396147261928e-14
+ k2 = 0.012897216193958 lk2 = 1.36104488355559e-08 wk2 = 3.14464223016169e-09 pk2 = -2.12137564846707e-15
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 103781.408935745 lvsat = -0.0308383331280536 wvsat = -0.228895417822604 pvsat = 1.54412848863129e-7
+ ua = -7.9435789278744e-09 lua = 6.94141918568807e-15 wua = 3.12788801261029e-14 pua = -2.1100732533069e-20
+ ub = 6.03901842708801e-18 lub = -4.26210824691357e-24 wub = -1.83388154951204e-23 pub = 1.23713649330082e-29
+ uc = 9.85959464678481e-12 luc = -8.31471122872103e-18 wuc = -3.74666853457179e-17 puc = 2.52750259342213e-23
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = -0.0158476594104472 lu0 = 2.29827176382877e-08 wu0 = 1.15366562464682e-07 pu0 = -7.78262830386744e-14
+ a0 = 1.06792881481362 la0 = -1.51392932473268e-07 wa0 = -6.82187415595184e-07 pa0 = 4.6020363056051e-13
+ keta = 0.20439965836152 lketa = -1.81865183530682e-07 wketa = -9.79383372029536e-07 pketa = 6.60692022771125e-13
+ a1 = 0.0
+ a2 = 0.5
+ ags = -2.44143323151152 lags = 2.13345840997767e-06 wags = 9.61351666293579e-06 pags = -6.48527834081649e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {0.124786874212527+0*(0.009/sqrt(l*w*mult))} lvoff = -1.33306495236371e-07 wvoff = -6.0068863177222e-07 pvoff = 4.05224550993539e-13
+ nfactor = {2.08600308605776+0*(0.02/sqrt(l*w*mult))} lnfactor = -1.80646469854565e-07 wnfactor = -2.31649251914335e-06 pnfactor = 1.56270585341411e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -0.138512393522682 leta0 = 9.39204857924018e-08 weta0 = 4.2660016546023e-07 peta0 = -2.87784471619471e-13
+ etab = -0.00179416616 letab = 8.51511259536e-10
+ dsub = 0.074039727213147 ldsub = 1.35448739868011e-07 wdsub = 6.10367058940381e-07 pdsub = -4.11753617961181e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.790310823914572 lpclm = 1.18899496250277e-06 wpclm = 5.35767965535723e-06 ppclm = -3.61429069550399e-12
+ pdiblc1 = -0.202026444642355 lpdiblc1 = 4.44550440881733e-07 wpdiblc1 = 2.00317618142681e-06 ppdiblc1 = -1.35134265199053e-12
+ pdiblc2 = 0.0473540801773804 lpdiblc2 = -2.42472518080608e-08 wpdiblc2 = -1.09259856295784e-07 ppdiblc2 = 7.3706699057136e-14
+ pdiblcb = -0.025
+ drout = -2.31616214999299 ldrout = 1.85377212949527e-06 wdrout = 8.35323021664869e-06 pdrout = -5.63508910415121e-12
+ pscbe1 = 475677157.72736 lpscbe1 = -51.0518106028774 wpscbe1 = -230.043121351 ppscbe1 = 0.000155187089663385
+ pscbe2 = 6.55695871368432e-09 lpscbe2 = 4.68621433074855e-15 wpscbe2 = 2.11164179925172e-14 ppscbe2 = -1.42451355777521e-20
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -0.000308907728446942 lalpha0 = 2.20019372966907e-10 walpha0 = 9.91423080147216e-10 palpha0 = -6.68814009867312e-16
+ alpha1 = 0.0
+ beta0 = 1.00632008888408 lbeta0 = 2.99120405260388e-05 wbeta0 = 0.00013478580068617 pbeta0 = -9.09265011428906e-11
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 5.95319590042466e-08 lagidl = -2.88903919442648e-14 wagidl = -9.40284381063768e-14 pagidl = 6.34315843465618e-20
+ bgidl = 2405869767.1954 lbgidl = -403.795164950017 wbgidl = -1819.52998404151 pbgidl = 0.0012274549272344
+ cgidl = 2254.11820666 lcgidl = -0.00116983614221284 wcgidl = -0.00527136558813224 pcgidl = 3.55606322575401e-9
+ egidl = -1.22811711014564 legidl = 1.15299534246625e-06 wegidl = 5.1954797362104e-06 pegidl = -3.50487063004754e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.790134844758 lkt1 = 1.00943666273747e-07 wkt1 = 4.90782313377829e-07 pkt1 = -3.31081748604683e-13
+ kt2 = -0.019032
+ at = 41611 lat = -0.0112057806
+ ute = -1.71258403862 lute = 1.57036112453052e-07 wute = 5.45313681530921e-07 pute = -3.67868609560759e-13
+ ua1 = 5.53349200000001e-10 lua1 = -6.40330320000131e-19
+ ub1 = -4.2831041e-18 lub1 = 4.6696088586e-25
+ uc1 = -2.69861592e-10 luc1 = 1.083823099632e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.02e-6
+ sbref = 2.01e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.47 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 6e-07 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.02/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.08790409285269+0*(0.0/sqrt(l*w*mult))} lvth0 = 2.6875486095109e-08 wvth0 = 1.21652637395119e-06 pvth0 = -3.53381275525226e-13
+ k1 = 0.353550686094241 lk1 = 9.72518223209012e-08 wk1 = 7.63631572736911e-07 pk1 = -3.36644384407245e-13
+ k2 = 0.081193984996048 lk2 = -1.8803197637916e-08 wk2 = -2.15269649772039e-07 pk2 = 1.01538047335777e-13
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 143181.725363993 lvsat = -0.0495377233049002 wvsat = -0.633750656679902 pvsat = 3.46557145224802e-7
+ ua = 1.97634927087013e-08 lua = -6.20835701303077e-15 wua = -5.5805025885567e-14 pua = 2.02292892600695e-20
+ ub = -1.62717155027567e-17 lub = 6.32656607619073e-24 wub = 4.42876382241169e-23 pub = -1.73511500021418e-29
+ uc = -1.48363103324958e-10 luc = 6.67777812286681e-17 wuc = 8.25354516886901e-16 puc = -3.8421991664538e-22
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0608632826600429 lu0 = -1.34242954683669e-08 wu0 = -1.55333192768222e-07 pu0 = 5.06478207948618e-14
+ a0 = 1.2847244170352 la0 = -2.54284125287631e-07 wa0 = -2.27778880591193e-06 pa0 = 1.21747605040484e-12
+ keta = -0.139656756606912 lketa = -1.85760089866634e-08 wketa = -1.85927898983486e-07 pketa = 2.8411805526347e-13
+ a1 = 0.0
+ a2 = 0.5
+ ags = -0.970108199456963 lags = 1.43516754976458e-06 wags = 1.11888924231904e-05 pags = -7.23295167663332e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.171361818960036+0*(0.009/sqrt(l*w*mult))} lvoff = 7.24567454332774e-09 wvoff = 8.4147565715014e-07 pvoff = -2.79226620529013e-13
+ nfactor = {7.70025551038833+0*(0.02/sqrt(l*w*mult))} lnfactor = -2.84517067044185e-06 wnfactor = -1.83648981403531e-05 pnfactor = 9.17927916124026e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 5.719768954e-05 lcit = -2.2400023455684e-11 wcit = -1.43471347872934e-10 pcit = 6.80915017004945e-17
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.719887544219851 leta0 = -3.13476124660204e-07 weta0 = -3.82228248661168e-06 peta0 = 1.72873523505386e-12
+ etab = 0.010539062546868 letab = -5.00183908474357e-09 wetab = 1.39999341254409e-07 petab = -6.64436873593425e-14
+ dsub = 0.632858182429997 ldsub = -1.29766498977906e-07 wdsub = -1.29708813450526e-06 pdsub = 4.93524616848119e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.409428155875322 lpclm = 6.19598842694485e-07 wpclm = 5.88433302672313e-06 ppclm = -3.86424038555425e-12
+ pdiblc1 = 0.857826518579751 lpdiblc1 = -5.84557754634792e-08 wpdiblc1 = 1.82890224624112e-06 ppdiblc1 = -1.2686322423514e-12
+ pdiblc2 = -0.0711581027940727 lpdiblc2 = 3.19986302301908e-08 wpdiblc2 = 3.37334344345194e-07 ppdiblc2 = -1.38246908567072e-13
+ pdiblcb = -1.1637075816 lpdiblcb = 5.4043061822736e-07 wpdiblcb = 5.73885391491736e-06 ppdiblcb = -2.72366006801978e-12
+ drout = 6.41712941042888 ldrout = -2.29104804508095e-06 wdrout = -2.46643839641092e-05 pdrout = 1.00350705860365e-11
+ pscbe1 = 846404983.179482 lpscbe1 = -226.999236562454 wpscbe1 = -996.540188873363 ppscbe1 = 0.000518966597909499
+ pscbe2 = 2.42949386975674e-08 lpscbe2 = -3.73223096960237e-15 wpscbe2 = -4.46406295335772e-14 ppscbe2 = 1.69631591781323e-20
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.000318009937487515 lalpha0 = -7.75157512855865e-11 walpha0 = -7.1796473753946e-10 palpha0 = 1.42461448406785e-16
+ alpha1 = 5.693537908e-10 lalpha1 = -2.7021530911368e-16 walpha1 = -2.86942695745868e-15 palpha1 = 1.36183003400989e-21
+ beta0 = -156.040962658619 lbeta0 = 0.000104446680918004 wbeta0 = 0.00109438292766258 pbeta0 = -5.46351297605895e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -2.33801581297652e-08 lagidl = 1.04596988475373e-14 wagidl = 5.41694143777317e-14 pagidl = -6.90311644239615e-21
+ bgidl = -1454027607.4344 lbgidl = 1428.11212904929 wbgidl = 16600.2615349239 pbgidl = -0.00751457812766657
+ cgidl = -401.103177254641 lcgidl = 9.03319265930526e-05 wcgidl = -2.88116204047728e-05 pcgidl = 1.06794711267055e-9
+ egidl = 10.7230360921119 legidl = -4.51902196732517e-06 wegidl = -4.84301351477103e-05 pegidl = 2.19458461938612e-11
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.588988457932 lkt1 = 5.47959108612712e-09 wkt1 = -8.09399009308137e-07 pkt1 = 2.85984307142076e-13
+ kt2 = -0.019032
+ at = 18000.0
+ ute = -0.847198531959997 lute = -2.53675849007785e-07 wute = -3.96005432052052e-06 pute = 1.77037904421286e-12
+ ua1 = 5.52e-10
+ ub1 = -4.8170792e-18 lub1 = 7.20385468320002e-25
+ uc1 = -4.1496e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 1.81e-6
+ sbref = 1.81e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.48 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 1.5e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.968873354504+0*(0.0/sqrt(l*w*mult))} wvth0 = 8.27260859638415e-8
+ k1 = 0.609396653813333 wk1 = -4.31245335151557e-8
+ k2 = 0.017373957190616 wk2 = 9.78237604755426e-9
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 220171.3276 wvsat = -0.0613167209531696
+ ua = 2.73094509798512e-09 wua = -7.87181255197357e-17
+ ub = -1.49470039626667e-19 wub = -6.82129017830172e-26
+ uc = -5.67301131333333e-11 wuc = 5.09412452702541e-17
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0203395130912 wu0 = -1.71874045297739e-9
+ a0 = 0.83004740837136 wa0 = 2.01038524502614e-7
+ keta = -0.00618613582613333 wketa = -5.2885281766632e-9
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.118208115626773 wags = 2.60807942185969e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0872410845777173+0*(0.009/sqrt(l*w*mult))} wvoff = -1.81280435949652e-8
+ nfactor = {1.93106812864+0*(0.02/sqrt(l*w*mult))} wnfactor = -3.54981688327357e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.51326533333333e-05 wcit = -1.56022190720533e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.080000000000001
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.69474425650536 wpclm = 2.36579877157297e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00463537189820613 wpdiblc2 = -5.15119026737021e-9
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 452172497.994453 wpscbe1 = -360.093224930867
+ pscbe2 = 1.501717205188e-08 wpscbe2 = -4.92874100486168e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 8.19931447648347e-05 walpha0 = -9.52245150301214e-11
+ alpha1 = 0.0
+ beta0 = 39.0839774229547 wbeta0 = -2.48634466777192e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.98819900666667e-08 wagidl = -1.55242079766931e-14
+ bgidl = 1758248978.66667 wbgidl = 53.0475448449806
+ cgidl = 1546.11431466667 wcgidl = -0.00166007610926647
+ egidl = 0.48984577703952 wegidl = 6.19092370655375e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.555469386666666 wkt1 = -6.24088762882132e-8
+ kt2 = -0.019032
+ at = 558874.883386667 wat = -0.334605190219256
+ ute = -1.51556938666667 wute = -6.24088762882132e-8
+ ua1 = 2.2096e-11
+ ub1 = -3.5693883624e-18 wub1 = -2.83648342729933e-25
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.49 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 1.5e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.968873354504+0*(0.0/sqrt(l*w*mult))} wvth0 = 8.27260859638411e-8
+ k1 = 0.609396653813333 wk1 = -4.31245335151553e-8
+ k2 = 0.017373957190616 wk2 = 9.78237604755423e-9
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 220171.3276 wvsat = -0.0613167209531698
+ ua = 2.73094509798512e-09 wua = -7.87181255197372e-17
+ ub = -1.49470039626667e-19 wub = -6.82129017830171e-26
+ uc = -5.67301131333333e-11 wuc = 5.09412452702541e-17
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0203395130912 wu0 = -1.71874045297739e-9
+ a0 = 0.83004740837136 wa0 = 2.01038524502614e-7
+ keta = -0.00618613582613333 wketa = -5.28852817666319e-9
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.118208115626773 wags = 2.60807942185968e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0872410845777173+0*(0.009/sqrt(l*w*mult))} wvoff = -1.81280435949651e-8
+ nfactor = {1.93106812864+0*(0.02/sqrt(l*w*mult))} wnfactor = -3.54981688327358e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.51326533333333e-05 wcit = -1.56022190720533e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.080000000000001
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.69474425650536 wpclm = 2.36579877157297e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00463537189820613 wpdiblc2 = -5.15119026737021e-9
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 452172497.994453 wpscbe1 = -360.093224930867
+ pscbe2 = 1.501717205188e-08 wpscbe2 = -4.92874100486042e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 8.19931447648347e-05 walpha0 = -9.52245150301214e-11
+ alpha1 = 0.0
+ beta0 = 39.0839774229547 wbeta0 = -2.48634466777189e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.98819900666667e-08 wagidl = -1.55242079766931e-14
+ bgidl = 1758248978.66667 wbgidl = 53.0475448449833
+ cgidl = 1546.11431466667 wcgidl = -0.00166007610926647
+ egidl = 0.48984577703952 wegidl = 6.19092370655375e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.555469386666667 wkt1 = -6.24088762882136e-8
+ kt2 = -0.019032
+ at = 558874.883386667 wat = -0.334605190219256
+ ute = -1.51556938666667 wute = -6.24088762882132e-8
+ ua1 = 2.2096e-11
+ ub1 = -3.5693883624e-18 wub1 = -2.83648342729933e-25
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.50 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 1.5e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.980311749270664+0*(0.0/sqrt(l*w*mult))} lvth0 = 9.00727834295713e-08 wvth0 = 1.00338880471971e-07 pvth0 = -1.38693711633721e-13
+ k1 = 0.627358094025273 lk1 = -1.41439157092943e-07 wk1 = -7.07814873077399e-08 pk1 = 2.17787448335085e-13
+ k2 = 0.0127182341077453 lk2 = 3.66619569883734e-08 wk2 = 1.69512398276661e-08 pk2 = -5.64519347228693e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 367572.917273724 lvsat = -1.16072855804471 wvsat = -0.288285099126411 pvsat = 1.78728519076301e-6
+ ua = 2.21945944214846e-09 lua = 4.02774494545134e-15 wua = 7.08865441394924e-16 pua = -6.20190555602619e-21
+ ub = 3.53587696232772e-19 lub = -3.96137844679874e-24 wub = -8.42819191228437e-25 pub = 6.09971468686691e-30
+ uc = -8.00367994323895e-11 luc = 1.83530831930548e-16 wuc = 8.68287876067956e-17 puc = -2.82600040883329e-22
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0189960366233255 lu0 = 1.05793397939246e-08 wu0 = 3.499392383499e-10 pu0 = -1.62900250973259e-14
+ a0 = 0.868206223096771 la0 = -3.00485402436721e-07 wa0 = 1.42281734223686e-07 pa0 = 4.62686220730452e-13
+ keta = -0.000222348776090169 lketa = -4.69624375042699e-08 wketa = -1.44715436211715e-08 pketa = 7.23125734193247e-14
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.0780716579990761 lags = 3.16058549235066e-07 wags = 8.78827511278947e-08 pags = -4.86665689877957e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0903981953872545+0*(0.009/sqrt(l*w*mult))} lvoff = 2.48609847807815e-08 wvoff = -1.3266736998883e-08 pvoff = -3.82808449215087e-14
+ nfactor = {1.91397040795738+0*(0.02/sqrt(l*w*mult))} lnfactor = 1.34637711287381e-07 wnfactor = -3.28654686411138e-07 pnfactor = -2.07314609289464e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.51326533333333e-05 wcit = -1.56022190720533e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.080000000000001
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -2.16471602210644 lpclm = 1.15754396654023e-05 wpclm = 4.62925541635845e-06 ppclm = -1.78238156950278e-11
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00787586638740351 lpdiblc2 = -2.55175979046336e-08 wpdiblc2 = -1.01408907198584e-08 ppdiblc2 = 3.92918951831632e-14
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 910950533.274049 lpscbe1 = -3612.6935166127 wpscbe1 = -1066.51780854225 ppscbe1 = 0.00556281102610617
+ pscbe2 = -4.58792987686793e-08 lpscbe2 = 4.79535349123576e-13 wpscbe2 = 9.37188547735653e-14 ppscbe2 = -7.38386612439086e-19
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.000137200722979547 lalpha0 = -4.34737595409577e-10 walpha0 = -1.80232923134823e-10 palpha0 = 6.69407210461286e-16
+ alpha1 = 0.0
+ beta0 = 40.8399525970386 lbeta0 = -1.38276021058414e-05 wbeta0 = -5.19018821692568e-06 pbeta0 = 2.12916864121663e-11
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 3.043310931685e-08 lagidl = -8.30858436474937e-14 wagidl = -3.17707791936484e-14 pagidl = 1.27935249705036e-19
+ bgidl = 1589234770.77071 lbgidl = 1330.91928149753 wbgidl = 313.294946106347 pbgidl = -0.00204934418597277
+ cgidl = 2213.53395095733 lcgidl = -0.00525566266793449 wcgidl = -0.0026877661955483 pcgidl = 8.09264835343485e-9
+ egidl = 1.52588651966067 legidl = -8.15840643184448e-06 wegidl = -9.76199020669694e-07 pegidl = 1.25622815901284e-11
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.555469386666667 wkt1 = -6.24088762882132e-8
+ kt2 = -0.019032
+ at = 989046.468965304 lat = -3.38742916779754 wat = -0.9969816770069 pat = 5.21594988285798e-6
+ ute = -1.47630940806133 lute = -3.09156627525558e-07 wute = -1.2286123430479e-07 pute = 4.76038138437343e-13
+ ua1 = 2.2096e-11
+ ub1 = -3.39095175963876e-18 lub1 = -1.40511687210366e-24 wub1 = -5.58404309915278e-25 pub1 = 2.16359333919772e-30
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.51 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 1.5e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.927648321915252+0*(0.0/sqrt(l*w*mult))} lvth0 = -1.13976932201711e-07 wvth0 = 9.8379505277999e-09 pvth0 = 2.11961191527964e-13
+ k1 = 0.623752670011104 lk1 = -1.27469581207642e-07 wk1 = -6.52298698324179e-08 pk1 = 1.96277151265202e-13
+ k2 = 0.0192934864694627 lk2 = 1.11854841876633e-08 wk2 = 9.76659440296284e-09 pk2 = -2.86143075603139e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 46535.1605493067 lvsat = 0.0831643341597204 wvsat = 0.20604755452682 pvsat = -1.28056109081801e-7
+ ua = 3.9585387692864e-09 lua = -2.71049181547732e-15 wua = -1.96849624204959e-15 pua = 4.17180002264792e-21
+ ub = -2.57219209403114e-18 lub = 7.37484792855782e-24 wub = 3.56892093304392e-24 pub = -1.09940135986388e-29
+ uc = -9.84849893595432e-11 luc = 2.55010188622297e-16 wuc = 1.33899355890493e-16 puc = -4.64979664755342e-22
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0205821450111916 lu0 = 4.43380423429879e-09 wu0 = -2.24213911242984e-09 pu0 = -6.2467583193947e-15
+ a0 = 0.602511664489173 la0 = 7.28974734344277e-07 wa0 = 6.89606600968494e-07 pa0 = -1.65797870795899e-12
+ keta = -0.000649818599090142 lketa = -4.53061629280742e-08 wketa = -1.38133272975954e-08 pketa = 6.97622484519969e-14
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.0877376435318664 lags = 2.78606721689717e-07 wags = 9.66510126330294e-08 pags = -5.20639195905752e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0292450521585447+0*(0.009/sqrt(l*w*mult))} lvoff = -2.12082983973178e-07 wvoff = -1.07430102329878e-07 pvoff = 3.26564530389963e-13
+ nfactor = {2.75513593974406+0*(0.02/sqrt(l*w*mult))} lnfactor = -3.1245422581733e-06 wnfactor = -1.49355246118491e-06 pnfactor = 4.30619830884898e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.51326533333333e-05 wcit = -1.56022190720533e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -0.0411860069686922 leta0 = 4.69547302600899e-07 weta0 = 1.86601728786366e-07 peta0 = -7.23007058355654e-13
+ etab = -0.174265553205729 letab = 4.03987312450918e-07 wetab = 1.60547681763969e-07 petab = -6.22058047762674e-13
+ dsub = 1.06687282068332 ldsub = -1.96392943101959e-06 wdsub = -7.80480741796893e-07 pdsub = 3.02405068216624e-12
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.25337585908138 lpclm = -1.66829913744805e-06 wpclm = -6.33908789927032e-07 ppclm = 2.56884033864596e-12
+ pdiblc1 = 0.77116114317852 lpdiblc1 = -1.47684696535949e-06 wpdiblc1 = -5.86910403621712e-07 ppdiblc1 = 2.27404304987269e-12
+ pdiblc2 = -0.00353185065671196 lpdiblc2 = 1.86827425544962e-08 wpdiblc2 = 7.42466635380245e-09 ppdiblc2 = -2.8767612254443e-14
+ pdiblcb = 0.354893438773333 lpdiblcb = -1.47193511787116e-06 wpdiblcb = -5.84958397449423e-07 ppdiblcb = 2.26647980675754e-12
+ drout = -0.275765565301332 ldrout = 3.23825725931654e-06 wdrout = 1.28690847438873e-06 pdrout = -4.98625557486658e-12
+ pscbe1 = -531169244.490317 lpscbe1 = 1974.94377431311 wpscbe1 = 1154.05245678021 ppscbe1 = -0.00304101052391223
+ pscbe2 = 1.37679714467424e-07 lpscbe2 = -2.3168240356103e-13 wpscbe2 = -1.88924579571334e-13 ppscbe2 = 3.5674363827366e-19
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 6.78184616996318e-05 lalpha0 = -1.65909085854416e-10 walpha0 = -7.33983947450542e-11 palpha0 = 2.55466146762286e-16
+ alpha1 = -1.89946719386667e-10 lalpha1 = 7.35967558935578e-16 walpha1 = 2.92479198724712e-16 palpha1 = -1.13323990337877e-21
+ beta0 = 102.55872450918 lbeta0 = -0.000252963155756623 wbeta0 = -0.000100224506332153 pbeta0 = 3.89511655381425e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.89666573427265e-08 lagidl = -3.86579288285547e-14 wagidl = -2.88359403758609e-14 pagidl = 1.16563923221637e-19
+ bgidl = 2966981482.86789 lbgidl = -4007.29812919423 wbgidl = -1531.19410343953 pbgidl = 0.0050973130853977
+ cgidl = 1925.05326817617 lcgidl = -0.0041379154144306 wcgidl = -0.0033000243729902 pcgidl = 1.04649038877512e-8
+ egidl = -4.06387392638522 legidl = 1.34996793924049e-05 wegidl = 7.63089175510998e-06 pegidl = -2.07867523297075e-11
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.551595850697333 lkt1 = -1.50084024667783e-08 wkt1 = -7.70328362244489e-08 pkt1 = 5.66619951689387e-14
+ kt2 = -0.019032
+ at = 176641.376237125 lat = -0.239684395512936 wat = 0.326220002250935 pat = 8.90726564055717e-8
+ ute = -1.61724830224533 lute = 2.36925211879769e-07 wute = -1.16991679489884e-07 pute = 4.5329596135151e-13
+ ua1 = -4.749579392e-10 lua1 = 1.92588519282432e-15 wua1 = -4.93038065763132e-32 pua1 = -3.29138418230241e-37
+ ub1 = -3.53462625911592e-18 lub1 = -8.48435656429458e-25 wub1 = 3.83440229528098e-25 pub1 = -1.48567751332956e-30
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.52 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 1.5e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.05362335866451+0*(0.0/sqrt(l*w*mult))} lvth0 = 1.22175871688446e-07 wvth0 = 2.02533434272605e-07 pvth0 = -1.49265762300047e-13
+ k1 = 0.536878287437307 lk1 = 3.53851363651982e-08 wk1 = 6.85389569571846e-08 pk1 = -5.44858914345865e-14
+ k2 = 0.0157659373009994 lk2 = 1.77982278588645e-08 wk2 = 8.38598213936976e-09 pk2 = -2.60262118109823e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 220505.293789662 lvsat = -0.242960077612651 wvsat = -0.0214297933081472 pvsat = 2.98372927169628e-7
+ ua = 4.19199147480626e-09 lua = -3.14812225724485e-15 wua = -2.32956028186381e-15 pua = 4.84865067168367e-21
+ ub = 1.32378817514904e-18 lub = 7.1443315952655e-26 wub = -2.19441657062925e-24 pub = -1.90061114253043e-31
+ uc = 7.01142326467686e-11 luc = -6.10459129507348e-17 wuc = -2.11576456718913e-16 puc = 1.8264929356225e-22
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0306356439247957 lu0 = -1.44124848291435e-08 wu0 = -1.70745871241426e-08 pu0 = 2.1558148723362e-14
+ a0 = 1.16602258977494 la0 = -3.27382846196429e-07 wa0 = -4.90056669864708e-07 pa0 = 5.53418059544935e-13
+ keta = 0.0949111547369622 lketa = -2.24444763543838e-07 wketa = -1.60957731796556e-07 pketa = 3.45599149125748e-13
+ a1 = 0.0
+ a2 = 0.5
+ ags = -0.722752703269909 lags = 1.79795192580432e-06 wags = 1.36753287564589e-06 pags = -2.90303433630966e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.217986347941804+0*(0.009/sqrt(l*w*mult))} lvoff = 1.4173144910212e-07 wvoff = 1.83192989952002e-07 pvoff = -2.18237518401649e-13
+ nfactor = {0.263168755464432+0*(0.02/sqrt(l*w*mult))} lnfactor = 1.54689942547729e-06 wnfactor = 2.10120096300197e-06 pnfactor = -2.43252646013174e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 2.39946719386667e-05 lcit = -1.66127400775579e-11 wcit = -2.92479198724712e-11 pcit = 2.55802307204633e-17
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.448611646210733 leta0 = -4.48627378049252e-07 weta0 = -5.67586738388701e-07 peta0 = 6.90794642210726e-13
+ etab = 0.0144628459367915 letab = 5.01970554183489e-08 wetab = -1.30055552322088e-07 petab = -7.72932251449519e-14
+ dsub = 0.00887034007083098 ldsub = 1.940201913658e-08 wdsub = 8.48627245840295e-07 pdsub = -2.9875151458429e-14
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.695449409891314 lpclm = 1.98496871176816e-06 wpclm = 2.36688758055655e-06 ppclm = -3.05645253746256e-12
+ pdiblc1 = -0.38920691316541 lpdiblc1 = 6.98378993062837e-07 wpdiblc1 = 1.19981968806445e-06 ppdiblc1 = -1.07536118000218e-12
+ pdiblc2 = 0.0105505347467062 lpdiblc2 = -7.7160971227516e-09 wpdiblc2 = -1.42593343608393e-08 ppdiblc2 = 1.18812154852244e-14
+ pdiblcb = -0.784786877546667 lpdiblcb = 6.64509603102315e-07 wpdiblcb = 1.16991679489885e-06 ppdiblcb = -1.02320922881853e-12
+ drout = 2.49616977591333 ldrout = -1.95801273132446e-06 wdrout = -2.98130647627224e-06 pdrout = 3.01494017164247e-12
+ pscbe1 = 644417705.399139 lpscbe1 = -228.811521949664 wpscbe1 = -656.111626311773 ppscbe1 = 0.000352323066252005
+ pscbe2 = 1.40691520276719e-08 lpscbe2 = 3.79567885291997e-17 wpscbe2 = 1.41047003114696e-15 ppscbe2 = -5.84457111501124e-23
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -0.000140877386537716 lalpha0 = 2.25312151251315e-10 walpha0 = 2.4795063758742e-10 palpha0 = -3.46934749248171e-16
+ alpha1 = 3.79893438773333e-10 lalpha1 = -3.32254801551158e-16 walpha1 = -5.84958397449424e-16 palpha1 = 5.11604614409266e-22
+ beta0 = -115.9577660173 lbeta0 = 0.000156667857384316 wbeta0 = 0.000236246311714559 pbeta0 = -2.41236540128941e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -2.80977251684966e-09 lagidl = 2.16416658620674e-15 wagidl = 4.5626700018835e-14 pagidl = -2.30237424622602e-20
+ bgidl = 204233490.406506 lbgidl = 1171.74925747388 wbgidl = 2174.26421400034 pbgidl = -0.00184893907647509
+ cgidl = -1642.68703795448 lcgidl = 0.00255017056344192 wcgidl = 0.00521750241321256 pcgidl = -5.50205182566445e-9
+ egidl = 5.30163325447747 legidl = -4.05690036884028e-06 wegidl = -6.79007873995367e-06 pegidl = 6.24679896033878e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.471097872551999 lkt1 = -1.65909912298021e-07 wkt1 = -1.69617964419921e-07 pkt1 = 2.3022207648417e-13
+ kt2 = -0.019032
+ at = 47253.4539598451 lat = 0.0028662035880529 wat = 0.755187475826846 pat = -7.15069769559831e-7
+ ute = -1.45430651503467 lute = -6.85254624253474e-08 wute = 4.29435477739219e-08 pute = 1.53481384322781e-13
+ ua1 = 5.524e-10
+ ub1 = -4.33384490176816e-18 lub1 = 6.49779611086435e-25 wub1 = -7.66880459056195e-25 pub1 = 6.70713649490546e-31
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.81e-6
+ sbref = 2.81e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.53 pmos
* DC IV MOS Parameters
+ lmin = 8.0e-07 lmax = 1e-06 wmin = 1.5e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.70229239882195+0*(0.0/sqrt(l*w*mult))} lvth0 = -1.85098185789854e-07 wvth0 = -5.59485066269065e-07 pvth0 = 5.17195618273699e-13
+ k1 = 0.582914710190694 lk1 = -4.87831897491381e-09 wk1 = 2.06604896996507e-08 pk1 = -1.26113839711472e-14
+ k2 = 0.0518473969198837 lk2 = -1.37586167238117e-08 wk2 = -1.10075803373536e-07 pk2 = 7.75804657986055e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -462157.780108221 lvsat = 0.354097046818438 wvsat = 1.44607153971751 pvsat = -9.85103738694609e-7
+ ua = -8.6941900061011e-09 lua = 8.12213206595672e-15 wua = 2.43055282410013e-14 pua = -1.84463977504142e-20
+ ub = 1.01362451031181e-17 lub = -7.63593151324905e-24 wub = -1.98153462942145e-23 pub = 1.52212040219946e-29
+ uc = 1.16911499258253e-11 luc = -9.94908480299773e-18 wuc = -1.80388276601953e-17 puc = 1.3381283187495e-23
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = -0.0111965332003222 lu0 = 2.21739372844845e-08 wu0 = 6.85200133668765e-08 pu0 = -5.33028888660833e-14
+ a0 = 0.452475147017018 la0 = 2.96685747239653e-07 wa0 = 1.12402218724165e-06 pa0 = -8.58255308880286e-13
+ keta = -0.485307462465598 lketa = 2.83014439061521e-07 wketa = 1.01809661222942e-06 pketa = -6.85601780159369e-13
+ a1 = 0.0
+ a2 = 0.5
+ ags = 3.44743236758265 lags = -1.84929193716333e-06 wags = -8.688788624982e-06 pags = 5.8922244481395e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0363439372263786+0*(0.009/sqrt(l*w*mult))} lvoff = -1.71330033095906e-08 wvoff = -1.76477643830165e-07 pvoff = 9.63304179042352e-14
+ nfactor = {2.8381746115144+0*(0.02/sqrt(l*w*mult))} lnfactor = -7.05200696224016e-07 wnfactor = -3.23458059985475e-06 pnfactor = 2.23414809474275e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -1.1865e-05 lcit = 1.4750129e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -0.262593379328194 leta0 = 1.73392537287094e-07 weta0 = 9.07579402469464e-07 peta0 = -5.99385664583826e-13
+ etab = 0.303690078252799 letab = -2.02761081965231e-07 wetab = -9.1770198599604e-07 petab = 6.11582345746287e-13
+ dsub = -0.824480742040193 ldsub = 7.48250875550881e-07 wdsub = 3.66289984762922e-06 pdsub = -2.49123796898302e-12
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 4.22927368356186 lpclm = -2.32219410576598e-06 wpclm = -6.83139168541464e-06 ppclm = 4.98836250855584e-12
+ pdiblc1 = 0.238800312090213 lpdiblc1 = 1.49123873854269e-07 wpdiblc1 = -1.00277919793656e-07 ppdiblc1 = 6.17041878305124e-14
+ pdiblc2 = -0.0475774277601603 lpdiblc2 = 4.31226188857538e-08 wpdiblc2 = 4.76485592842999e-08 ppdiblc2 = -4.22634282968143e-14
+ pdiblcb = -0.025
+ drout = 0.0650139206247555 ldrout = 1.68276179710929e-07 wdrout = 8.34378872444574e-07 pdrout = -3.22258234345252e-13
+ pscbe1 = 217166683.079076 lpscbe1 = 144.862222171462 wpscbe1 = -780.435191960833 ppscbe1 = 0.000461056456768674
+ pscbe2 = 1.60998186969081e-08 lpscbe2 = -1.73806428038484e-15 wpscbe2 = 6.07843123897767e-15 ppscbe2 = -4.14104458351883e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.000505036354149857 lalpha0 = -3.39604006354036e-10 walpha0 = -8.10532718893197e-10 palpha0 = 5.78814794329778e-16
+ alpha1 = 0.0
+ beta0 = 130.575706723585 lbeta0 = -5.89503178748624e-05 wbeta0 = -0.000195189818262158 pbeta0 = 1.36097499148696e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -8.88076773265675e-08 lagidl = 7.7377934132786e-14 wagidl = 1.78616317101418e-13 pagidl = -1.39336461562687e-19
+ bgidl = 591087916.463999 lbgidl = 833.406376443998 wbgidl = 460.184331086402 pbgidl = -0.000349804810878549
+ cgidl = 3778.797520848 lcgidl = -0.00219145983168673 wcgidl = -0.00458886850548367 pcgidl = 3.07460017982727e-9
+ egidl = 0.172745124172152 legidl = 4.28825189924754e-07 wegidl = 4.89769816642074e-06 pegidl = -3.97533072197628e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.72925405816 lkt1 = 5.98734876347365e-08 wkt1 = 4.09371024012536e-07 pkt1 = -2.76161692798857e-13
+ kt2 = -0.019032
+ at = 119332.932413333 lat = -0.060174508267368 wat = -0.220287731078321 pat = 1.38080846399428e-7
+ ute = -1.71094430237333 lute = 1.55929946381049e-07 wute = 9.55199056029249e-07 pute = -6.44377283197332e-13
+ ua1 = 5.524e-10
+ ub1 = -3.5909e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.41e-6
+ sbref = 2.41e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.54 pmos
* DC IV MOS Parameters
+ lmin = 6e-07 lmax = 8.0e-07 wmin = 1.5e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.14070505548078+0*(0.0/sqrt(l*w*mult))} lvth0 = 1.10654992392189e-07 wvth0 = 4.71410935903689e-07 pvth0 = -1.78246824792042e-13
+ k1 = 0.698431172616079 lk1 = -8.28057245270793e-08 wk1 = -3.71162656113668e-07 pk1 = 2.51712510194518e-13
+ k2 = -0.019269157326313 lk2 = 3.42166107706726e-08 wk2 = 1.00923855791587e-07 pk2 = -6.4759904274187e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 30533.8222030737 lvsat = 0.0217272918992389 wvsat = -0.0062376966629768 pvsat = -5.3759278323346e-9
+ ua = 2.92985860259923e-09 lua = 2.80548874527483e-16 wua = -1.77415178528069e-15 pua = -8.53045604684336e-22
+ ub = -5.88810952315307e-19 lub = -4.00808698253699e-25 wub = 1.8084337410723e-24 pub = 6.33802010190126e-31
+ uc = -5.16175324670252e-12 luc = 1.41988367718952e-18 wuc = 8.19514789551333e-18 puc = -4.316156722386e-24
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0266087270777768 lu0 = -3.32949129912104e-09 wu0 = -1.36921913566756e-08 pu0 = 2.15746444042495e-15
+ a0 = 1.00432424117867 la0 = -7.55916516817951e-08 wa0 = -4.88842487077947e-07 pa0 = 2.29783200415714e-13
+ keta = -0.140377313152704 lketa = 5.03245603350429e-08 wketa = 6.8668286871517e-08 pketa = -4.51174318729289e-14
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.673145394727268 lags = 2.22420547249156e-08 wags = 1.4583301320963e-07 pags = -6.761130898458e-14
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0528562723687987+0*(0.009/sqrt(l*w*mult))} lvoff = -5.99378202251413e-09 wvoff = -6.06897053668912e-08 pvoff = 1.82198746169104e-14
+ nfactor = {0.929469309719281+0*(0.02/sqrt(l*w*mult))} lnfactor = 5.82411900366975e-07 wnfactor = 1.19913422803525e-06 pnfactor = -7.56835928151845e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.0236218310374699 leta0 = -1.9688243625583e-08 weta0 = -6.62548018208209e-08 peta0 = 5.75628896304012e-14
+ etab = 0.0105412241205351 letab = -5.00286496760594e-09 wetab = -3.74970700332094e-08 petab = 1.77961094377612e-14
+ dsub = 0.300823787619908 ldsub = -1.08795601578229e-08 wdsub = -7.90102207478494e-08 pdsub = 3.30545631441489e-14
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.658295427465204 lpclm = 8.67878257968195e-08 wpclm = 9.54212166837996e-07 ppclm = -2.63805850173789e-13
+ pdiblc1 = 0.324468714115882 lpdiblc1 = 9.13319698477532e-08 wpdiblc1 = 4.02738303814159e-07 ppdiblc1 = -2.77630556615321e-13
+ pdiblc2 = 0.0193771759787055 lpdiblc2 = -2.044956796485e-09 wpdiblc2 = -2.42157748202691e-08 ppdiblc2 = 6.21625149012792e-15
+ pdiblcb = -0.025
+ drout = 0.548770446357115 ldrout = -1.58065972548121e-07 wdrout = -3.55580430005974e-07 pdrout = 4.80488311087888e-13
+ pscbe1 = 357852922.138685 lpscbe1 = 49.9552853018504 wpscbe1 = 128.118518694513 ppscbe1 = -0.000151853876439423
+ pscbe2 = 1.62782400568239e-08 lpscbe2 = -1.85842732978404e-15 wpscbe2 = -8.43429414923316e-15 ppscbe2 = 5.64923996336819e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -5.20084508724032e-06 lalpha0 = 4.60200825131024e-12 walpha0 = 6.82161109379287e-11 palpha0 = -1.39891662742999e-17
+ alpha1 = 0.0
+ beta0 = 44.9622091207737 lbeta0 = -1.19545239200562e-06 wbeta0 = 1.16886503058862e-06 pbeta0 = 3.63393139940911e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.45595420486649e-07 lagidl = -8.07503956520101e-14 wagidl = -3.55643804066739e-13 pagidl = 2.21075416177352e-19
+ bgidl = 1242353569.64107 lbgidl = 394.06256681075 wbgidl = 1717.32189921936 pbgidl = -0.00119786981434105
+ cgidl = 1641.06182269866 lcgidl = -0.000749343329715186 wcgidl = -0.00340779924439211 pcgidl = 2.2778508562949e-9
+ egidl = 3.36880945771576 legidl = -1.72723980948376e-06 wegidl = -8.77823925706842e-06 pegidl = 5.25045666390951e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.648170118176 lkt1 = 5.17426172152944e-09 wkt1 = 5.92385053727712e-08 pkt1 = -3.99622957244713e-14
+ kt2 = -0.019032
+ at = 39435.7815173334 lat = -0.00627589027292641 wat = 0.00661222044273618 pat = -1.4985860896677e-8
+ ute = -1.2503778607208 lute = -1.54768175157749e-07 wute = -8.59698809222354e-07 pute = 5.79952816701402e-13
+ ua1 = 5.533492e-10 lua1 = -6.40330320000131e-19
+ ub1 = -8.00659583948808e-19 lub1 = -1.88229618466814e-24 wub1 = -1.05859209101144e-23 pub1 = 7.14126224596315e-30
+ uc1 = -4.34785643143487e-10 luc1 = 2.19640074864597e-16 wuc1 = 5.01335470969769e-16 puc1 = -3.38200908716207e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.02e-6
+ sbref = 2.01e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.55 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 6e-07 wmin = 1.5e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.014/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.629115353200026+0*(0.0/sqrt(l*w*mult))} lvth0 = -1.32145480310255e-07 wvth0 = -1.78097801690021e-07 pvth0 = 1.30010022069931e-13
+ k1 = 0.440257151523626 lk1 = 3.97236658833982e-08 wk1 = 5.00061605950527e-07 pk1 = -1.61770524581149e-13
+ k2 = 0.0657381702874795 lk2 = -6.12786691483331e-09 wk2 = -1.68287126044191e-07 pk2 = 6.30076277050735e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -166485.425378911 lvsat = 0.115232626801649 wvsat = 0.307574309479776 pvsat = -1.54311105947685e-7
+ ua = 3.86166670608035e-09 lua = -1.61687251384656e-16 wua = -7.46671881010385e-15 pua = 1.84864670529673e-21
+ ub = -6.15810599683067e-18 lub = 2.24237872987329e-24 wub = 1.3544328502441e-23 pub = -4.93605364355547e-30
+ uc = 2.48879185694008e-10 luc = -1.19147945944071e-16 wuc = -3.82181004303794e-16 puc = 1.80956365111405e-22
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.00905916996511358 lu0 = 4.99952850654893e-09 wu0 = 2.14074178537311e-09 pu0 = -5.35684562879141e-15
+ a0 = 0.118525076307357 la0 = 3.44808631966128e-07 wa0 = 1.2672192852352e-06 pa0 = -6.03643716724102e-13
+ keta = -0.341161784217488 lketa = 1.45616870302389e-07 wketa = 4.26606277927031e-07 pketa = -2.14994802427876e-13
+ a1 = 0.0
+ a2 = 0.5
+ ags = 5.22923093699619 lags = -2.14007614363592e-06 wags = -7.65583388644335e-06 pags = 3.63505980159072e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {0.250812582547504+0*(0.009/sqrt(l*w*mult))} lvoff = -1.50115020565792e-07 wvoff = -4.41848399854877e-07 pvoff = 1.99117791020908e-13
+ nfactor = {2.29932446318389+0*(0.02/sqrt(l*w*mult))} lnfactor = -6.77213554673308e-08 wnfactor = -1.94716954678527e-06 pnfactor = 7.36399843377975e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -0.948417572241565 leta0 = 4.41641657170647e-07 weta0 = 1.24902473318727e-06 peta0 = -5.66668777684437e-13
+ etab = 0.0609898417717921 letab = -2.89457789048925e-08 wetab = -1.33607356303983e-08 petab = 6.34100513018702e-15
+ dsub = 0.145712301180307 ldsub = 6.27363513064119e-08 wdsub = 1.83735966734028e-07 pdsub = -9.16447774347503e-14
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 3.37409536909603 lpclm = -1.20213082650117e-06 wpclm = -3.12765050935632e-06 ppclm = 1.67344617594803e-12
+ pdiblc1 = 1.73500582942244 lpdiblc1 = -5.78108945076741e-07 wpdiblc1 = -8.37543914141252e-07 ppdiblc1 = 3.11007384026317e-13
+ pdiblc2 = 0.0573829501181448 lpdiblc2 = -2.00824972030629e-08 wpdiblc2 = -5.34042341331533e-08 ppdiblc2 = 2.00690942800228e-14
+ pdiblcb = 1.49327677546667 lpdiblcb = -7.20574157636481e-07 wpdiblcb = -2.33783650575648e-06 ppdiblcb = 1.10953720563202e-12
+ drout = -2.72219518707034 ldrout = 1.39433431707655e-06 wdrout = 3.11729839007053e-06 pdrout = -1.16773997692042e-12
+ pscbe1 = 713259447.622577 lpscbe1 = -118.720651692805 wpscbe1 = -591.804922469626 ppscbe1 = 0.000189821788737078
+ pscbe2 = 4.99114238570167e-09 lpscbe2 = 3.49842922493058e-15 wpscbe2 = 1.4038973280047e-14 ppscbe2 = -5.01657275856818e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 9.12820341035211e-05 lalpha0 = -4.11887662126251e-11 walpha0 = -2.8758163744408e-11 palpha0 = 3.20348244899371e-17
+ alpha1 = -7.59138387733334e-10 lalpha1 = 3.60287078818241e-16 walpha1 = 1.16891825287824e-15 palpha1 = -5.54768602816012e-22
+ beta0 = 355.409532267051 lbeta0 = -0.000148533751957229 wbeta0 = -0.000460322241010489 pbeta0 = 2.22657610326505e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -2.07668402267066e-07 lagidl = 8.69086146269033e-14 wagidl = 6.14368081753324e-13 pagidl = -2.3929222483285e-19
+ bgidl = 7062135380.33868 lbgidl = -2368.00588054633 wbgidl = -9287.13665065678 pbgidl = 0.00402484621343016
+ cgidl = -3615.63314697782 lcgidl = 0.00174548410289327 wcgidl = 0.00974270372343987 pcgidl = -3.96337785223815e-9
+ egidl = -13.9974850597707 legidl = 6.51480356851532e-06 wegidl = 2.67152061676978e-05 pegidl = -1.15947325346845e-11
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.985477574250668 lkt1 = 1.65260380374567e-07 wkt1 = 3.95847020520883e-07 pkt1 = -1.99716697013765e-13
+ kt2 = -0.019032
+ at = 6985.32594666662 lat = 0.00912509594091201 wat = 0.0334823621286266 pat = -2.77384301408006e-8
+ ute = -2.82015912002187 lute = 5.90250010506539e-07 wute = 2.03734338322759e-06 pute = -7.94983407835346e-13
+ ua1 = 5.52e-10
+ ub1 = -8.95945646613974e-18 lub1 = 1.98986881561968e-24 wub1 = 1.25919818441025e-23 pub1 = -3.85897040118818e-30
+ uc1 = 2.80042322559999e-11 wuc1 = -2.1126652801086e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 1.81e-6
+ sbref = 1.81e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.56 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 1e-06 wmax = 1.5e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.923308319008+0*(0.0/sqrt(l*w*mult))} wvth0 = 1.25652265672422e-8
+ k1 = 0.57419461168 wk1 = 1.10794301535827e-8
+ k2 = 0.02360999315408 wk2 = 1.8015281515624e-10
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 388712.640848 wvsat = -0.320835960927187
+ ua = 3.57135481382944e-09 wua = -1.37277764433796e-15
+ ub = -8.9425976928e-19 wub = 1.07861134477827e-24
+ uc = 2.0984334234544e-11 wuc = -6.87231499290139e-17
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.021507731812 wu0 = -3.51755896639035e-9
+ a0 = 1.0701681373768 wa0 = -1.68698413537048e-7
+ keta = -0.0126128169696 wketa = 4.6072497413222e-9
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.17292289325152 wags = -5.81688015088774e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.080992296419832+0*(0.009/sqrt(l*w*mult))} wvoff = -2.77499026053243e-8
+ nfactor = {1.67041750784+0*(0.02/sqrt(l*w*mult))} wnfactor = 4.6367094977999e-8
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 5.0e-6
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.080000000000001
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.41835776951608 wpclm = -2.42774327568674e-6
+ pdiblc1 = 0.39
+ pdiblc2 = -0.0031771021168272 wpdiblc2 = 6.87842597108206e-9
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 204999413.56688 wpscbe1 = 20.5029017783725
+ pscbe2 = 1.495696373248e-08 wpscbe2 = 4.34211193302208e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -7.1542079670088e-05 walpha0 = 1.41188409413875e-10
+ alpha1 = 0.0
+ beta0 = 34.203828731392 wbeta0 = 5.02808876690154e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -1.14118384e-08 wagidl = 3.26619039209664e-14
+ bgidl = 2358972901.6 wbgidl = -871.944748792073
+ cgidl = -1470.179744 wcgidl = 0.00298440141709223
+ egidl = -0.41413520492296 wegidl = 2.01103867075727e-6
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.67918368 wkt1 = 1.2808589772928e-7
+ kt2 = -0.019032
+ at = 737690.68416 wat = -0.609945044986832
+ ute = -1.5561
+ ua1 = 2.2096e-11
+ ub1 = -5.1612758248e-18 wub1 = 2.16753360432374e-24
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.57 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 1e-06 wmax = 1.5e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.923308319008+0*(0.0/sqrt(l*w*mult))} wvth0 = 1.25652265672431e-8
+ k1 = 0.57419461168 wk1 = 1.10794301535827e-8
+ k2 = 0.02360999315408 wk2 = 1.80152815156227e-10
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 388712.640848 wvsat = -0.320835960927187
+ ua = 3.57135481382944e-09 wua = -1.37277764433796e-15
+ ub = -8.9425976928e-19 wub = 1.07861134477827e-24
+ uc = 2.0984334234544e-11 wuc = -6.87231499290139e-17
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.021507731812 wu0 = -3.51755896639036e-9
+ a0 = 1.0701681373768 wa0 = -1.68698413537048e-7
+ keta = -0.0126128169696 wketa = 4.6072497413222e-9
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.17292289325152 wags = -5.81688015088775e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.080992296419832+0*(0.009/sqrt(l*w*mult))} wvoff = -2.77499026053243e-8
+ nfactor = {1.67041750784+0*(0.02/sqrt(l*w*mult))} wnfactor = 4.63670949780007e-8
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 5.0e-6
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.080000000000001
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.41835776951608 wpclm = -2.42774327568674e-6
+ pdiblc1 = 0.39
+ pdiblc2 = -0.0031771021168272 wpdiblc2 = 6.87842597108206e-9
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 204999413.56688 wpscbe1 = 20.5029017783727
+ pscbe2 = 1.495696373248e-08 wpscbe2 = 4.34211193302208e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -7.1542079670088e-05 walpha0 = 1.41188409413875e-10
+ alpha1 = 0.0
+ beta0 = 34.203828731392 wbeta0 = 5.02808876690154e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -1.14118384e-08 wagidl = 3.26619039209664e-14
+ bgidl = 2358972901.6 wbgidl = -871.944748792073
+ cgidl = -1470.179744 wcgidl = 0.00298440141709223
+ egidl = -0.41413520492296 wegidl = 2.01103867075727e-6
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.67918368 wkt1 = 1.2808589772928e-7
+ kt2 = -0.019032
+ at = 737690.68416 wat = -0.609945044986832
+ ute = -1.5561
+ ua1 = 2.2096e-11
+ ub1 = -5.1612758248e-18 wub1 = 2.16753360432375e-24
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.58 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 1e-06 wmax = 1.5e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.888906450614717+0*(0.0/sqrt(l*w*mult))} lvth0 = -2.70900952849742e-07 wvth0 = -4.04066327772603e-08 pvth0 = 4.17132203594222e-13
+ k1 = 0.6149861466937 lk1 = -3.21217021618882e-07 wk1 = -5.17312122943728e-08 pk1 = 4.94608685020668e-13
+ k2 = 0.0115917312511577 lk2 = 9.46390051807521e-08 wk2 = 1.86858244202284e-08 pk2 = -1.45724761621301e-13
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 469437.577842519 lvsat = -0.635676588857042 wvsat = -0.4451358960116 pvsat = 9.78812268815718e-7
+ ua = 2.99919982741506e-09 lua = 4.50549165601868e-15 wua = -4.91775684877037e-16 pua = -6.93753802997094e-21
+ ub = -6.29709038744236e-19 lub = -2.08323118267693e-24 wub = 6.71257188102219e-25 pub = 3.20775104216121e-30
+ uc = 5.16162993217801e-11 luc = -2.41214472275949e-16 wuc = -1.1589012724248e-16 puc = 3.71421079552617e-22
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0200867763157697 lu0 = 1.11894561506152e-08 wu0 = -1.32957737711688e-09 pu0 = -1.72294798228927e-14
+ a0 = 0.995145554817677 la0 = 5.90772828620065e-07 wa0 = -5.31789410028404e-08 pa0 = -9.09669638417864e-13
+ keta = -0.0159271040095032 lketa = 2.60986847244221e-08 wketa = 9.71057566821705e-09 pketa = -4.01866503439262e-14
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.161431384023011 lags = 9.04910385708161e-08 wags = -4.04742215648566e-08 pags = -1.39337739227188e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0596202535227175+0*(0.009/sqrt(l*w*mult))} lvoff = -1.68296288997617e-07 wvoff = -6.06584887701296e-08 pvoff = 2.59141952613376e-13
+ nfactor = {1.78630575521473+0*(0.02/sqrt(l*w*mult))} lnfactor = -9.12573592777009e-07 wnfactor = -1.32077164776613e-07 pnfactor = 1.40517716786366e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.5071983954e-05 lcit = -7.93128448441685e-11 wcit = -1.55088006044334e-11 pcit = 1.22125601239671e-16
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.080000000000001
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 4.09049065771566 lpclm = -1.31673776414164e-05 wpclm = -5.0024868084049e-06 ppclm = 2.02750754227424e-11
+ pdiblc1 = 0.39
+ pdiblc2 = -0.00750416058229188 lpdiblc2 = 3.40738545921481e-08 wpdiblc2 = 1.35412132879707e-08 ppdiblc2 = -5.24667850055713e-14
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 205686443.73635 lpscbe1 = -5.41008777251045 wpscbe1 = 19.445015471543 ppscbe1 = 8.33043151176032e-6
+ pscbe2 = 1.49744204950691e-08 lpscbe2 = -1.37465022683962e-16 wpscbe2 = 1.6541266122612e-17 ppscbe2 = 2.11668092068677e-22
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -0.000200952048093326 lalpha0 = 1.01905173734563e-09 walpha0 = 3.40453361152103e-10 palpha0 = -1.56913178895785e-15
+ alpha1 = 2.0143967908e-10 lalpha1 = -1.58625689688337e-15 walpha1 = -3.10176012088668e-16 palpha1 = 2.44251202479343e-21
+ beta0 = -38.3939800939154 lbeta0 = 0.000571678705375765 wbeta0 = 0.000116813904404874 pbeta0 = -8.80268583822781e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.59839579548801e-08 lagidl = -2.15730937976138e-13 wagidl = -9.52203372309247e-15 pagidl = 3.32181635371906e-19
+ bgidl = 2262080415.96252 lbgidl = 762.989567400902 wbgidl = -722.750086977425 pbgidl = -0.00117484828392564
+ cgidl = -3299.2520300464 lcgidl = 0.014403212623701 wcgidl = 0.00580079960685733 pcgidl = -2.21780091851243e-8
+ egidl = 0.552905787573086 legidl = -7.61506099950936e-06 wegidl = 5.21992818675833e-07 pegidl = 1.17256404668005e-11
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.719471615816 lkt1 = 3.17251379376672e-07 wkt1 = 1.90121100147013e-07 pkt1 = -4.88502404958682e-13
+ kt2 = -0.019032
+ at = 875797.728137248 lat = -1.08753772850324 wat = -0.822601718874822 pat = 1.67458624419837e-6
+ ute = -1.26260238758044 lute = -2.31117629875907e-06 wute = -4.5192644961319e-07 pute = 3.55874002012402e-12
+ ua1 = 2.2096e-11
+ ub1 = -3.79773063710748e-18 lub1 = -1.07373729350035e-23 wub1 = 6.79521784955446e-26 pub1 = 1.65333638958267e-29
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.59 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 1e-06 wmax = 1.5e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.949284647685332+0*(0.0/sqrt(l*w*mult))} lvth0 = -3.69595904799331e-08 wvth0 = 4.31534784032697e-08 pvth0 = 9.33701968141383e-14
+ k1 = 0.509433151301808 lk1 = 8.77586143265425e-08 wk1 = 1.10798867798081e-07 pk1 = -1.35130363305552e-13
+ k2 = 0.0546813629612557 lk2 = -7.23160818431938e-08 wk2 = -4.47235162675941e-08 pk2 = 9.99610698077358e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 112084.445402218 lvsat = 0.748923858096152 wvsat = 0.105115027907447 pvsat = -1.15318996100102e-6
+ ua = 3.54839045830371e-09 lua = 2.37759763757749e-15 wua = -1.33695151339169e-15 pua = -3.66281976480805e-21
+ ub = -9.84473278034896e-19 lub = -7.08661661121336e-25 wub = 1.12415785104817e-24 pub = 1.45294213351083e-30
+ uc = 6.09649992896399e-11 luc = -2.77436945171419e-16 wuc = -1.11621098831565e-16 puc = 3.54880302071687e-22
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0210188494257602 lu0 = 7.57804567864602e-09 wu0 = -2.914574823165e-09 pu0 = -1.10882487184348e-14
+ a0 = 1.55308049189583 la0 = -1.57100187858296e-06 wa0 = -7.74075477196975e-07 pa0 = 1.88351608071993e-12
+ keta = -0.213960348163508 lketa = 7.93398292523531e-07 wketa = 3.14641372883578e-07 pketa = -1.22167151723456e-12
+ a1 = 0.0
+ a2 = 0.5
+ ags = 1.34851015546059 lags = -4.50896436924121e-06 wags = -1.84468145814477e-06 pags = 6.85124361962533e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0817846755804622+0*(0.009/sqrt(l*w*mult))} lvoff = -8.24180192926798e-08 wvoff = -2.65298003433027e-08 pvoff = 1.26906936434791e-13
+ nfactor = {1.89978698059241+0*(0.02/sqrt(l*w*mult))} lnfactor = -1.35226794862538e-06 wnfactor = -1.76489555279027e-07 pnfactor = 1.57725741610432e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -1.13508613939187e-05 lcit = 2.30651117408773e-11 wcit = 2.51769909709104e-11 pcit = -3.55155667981559e-17
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -0.075936126527999 leta0 = 6.04190115845389e-07 weta0 = 2.40109823883308e-07 peta0 = -9.30329523618267e-13
+ etab = 0.0651810280871232 letab = -5.23772411426368e-07 wetab = -2.0815120632444e-07 petab = 8.06502664024675e-13
+ dsub = -0.0247604744799998 ldsub = 2.26571293442021e-06 wdsub = 9.00411839562406e-07 pdsub = -3.4887357135685e-12
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.62164579129454 lpclm = -7.47619132198113e-06 wpclm = -2.74076535846913e-06 ppclm = 1.15118094928213e-11
+ pdiblc1 = 0.391770459796567 lpdiblc1 = -6.85982352777981e-09 wpdiblc1 = -2.72614691291493e-09 ppdiblc1 = 1.0562728828781e-14
+ pdiblc2 = 0.00129
+ pdiblcb = -0.025
+ drout = 0.712038054729069 ldrout = -5.89086646853249e-07 wdrout = -2.34107588519601e-07 pdrout = 9.07073262478047e-13
+ pscbe1 = 369667836.56033 lpscbe1 = -640.772392408302 wpscbe1 = -233.05287727325 ppscbe1 = 0.000986658766740734
+ pscbe2 = 1.44721510918496e-08 lpscbe2 = 1.80862800703029e-15 wpscbe2 = 7.89933684122374e-16 ppscbe2 = -2.78491817071321e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.00068534710206513 lalpha0 = -2.41500294985833e-09 walpha0 = -1.02426652506529e-09 palpha0 = 3.71861188218005e-15
+ alpha1 = -4.0287935816e-10 lalpha1 = 7.55237644806736e-16 walpha1 = 6.20352024177336e-16 palpha1 = -1.16291190452283e-21
+ beta0 = 211.179349818911 lbeta0 = -0.000395318118704472 wbeta0 = -0.000267478110701576 pbeta0 = 6.08709257908671e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -5.666171561008e-08 lagidl = 6.5741988818656e-14 wagidl = 8.76163257833788e-14 pagidl = -4.41906523718677e-20
+ bgidl = 3272749501.13632 lbgidl = -3152.94887001351 wbgidl = -2002.01447489718 pbgidl = 0.00378178951350825
+ cgidl = -1016.5072153344 lcgidl = 0.00555848956461787 wcgidl = 0.00122937869327745 pcgidl = -4.46558171336768e-9
+ egidl = -2.47075335750202 legidl = 4.10040872399863e-06 wegidl = 5.17781107562589e-06 pegidl = -6.3137929515782e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.730929711172 lkt1 = 3.61646915643031e-07 wkt1 = 1.99104724799001e-07 pkt1 = -5.23310357035276e-13
+ kt2 = -0.019032
+ at = 344315.62126009 lat = 0.971742842803001 wat = 0.0680358704615553 pat = -1.77627815944436e-6
+ ute = -2.26852700534952 lute = 1.58637922524901e-06 wute = 8.8584466243513e-07 pute = -1.6245879306184e-12
+ ua1 = -4.42623577296637e-11 lua1 = 2.57112092859355e-16 wua1 = -6.63183333565698e-16 pua1 = 2.56957014423365e-21
+ ub1 = -5.90954616428688e-18 lub1 = -2.55493249339422e-24 wub1 = 4.04033239983072e-24 pub1 = 1.14197949024143e-30
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.60 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 1e-06 wmax = 1.5e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.968336646847426+0*(0.0/sqrt(l*w*mult))} lvth0 = -1.24471285067569e-09 wvth0 = 7.120929656351e-08 pvth0 = 4.07767600909523e-14
+ k1 = 0.561322215865327 lk1 = -9.51262610423199e-09 wk1 = 3.09002937394315e-08 pk1 = 1.46475036247914e-14
+ k2 = 0.0147381122176309 lk2 = 2.56153600080531e-09 wk2 = 9.96862309144029e-09 pk2 = -2.56481463471016e-15
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 637573.698695562 lvsat = -0.236158296127551 wvsat = -0.663630054908631 pvsat = 2.87899571245998e-7
+ ua = 3.51316879949182e-09 lua = 2.44362415918626e-15 wua = -1.28431184170534e-15 pua = -3.76149809335128e-21
+ ub = -1.77263632747885e-19 lub = -2.22185686217636e-24 wub = 1.168969989632e-25 pub = 3.34115332682931e-30
+ uc = -1.63252202640391e-10 luc = 1.42880621566616e-16 wuc = 1.47760246870513e-16 puc = -1.31355968581429e-22
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0218816507067476 lu0 = 5.96063839730704e-09 wu0 = -3.59522338296498e-09 pu0 = -9.81230492823374e-15
+ a0 = 0.502642764795155 la0 = 3.98148684639971e-07 wa0 = 5.31412931119872e-07 pa0 = -5.63752489510832e-13
+ keta = 0.259194789390787 lketa = -9.3578328335752e-08 wketa = -4.13921015301977e-07 pketa = 1.44091535658078e-13
+ a1 = 0.0
+ a2 = 0.5
+ ags = -0.962060637324138 lags = -1.77568361086969e-07 wags = 1.73601827527086e-06 pags = 1.38863899364403e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.113904474791415+0*(0.009/sqrt(l*w*mult))} lvoff = -2.22062436918282e-08 wvoff = 2.29281380025252e-08 pvoff = 3.41930852117024e-14
+ nfactor = {1.2387013094552+0*(0.02/sqrt(l*w*mult))} lnfactor = -1.12996749511567e-07 wnfactor = 5.99079838497198e-07 pnfactor = 1.23375030531401e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -2.58621302816268e-06 lcit = 6.63490191443108e-12 wcit = 1.16812204759128e-11 pcit = -1.02163954282333e-17
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.318286791015256 leta0 = -1.34820165381196e-07 weta0 = -3.66913047658125e-07 peta0 = 2.07595551373304e-13
+ etab = -0.214475151334308 letab = 4.71062517046849e-10 wetab = 2.22462260123962e-07 petab = -7.25340179498641e-16
+ dsub = 1.27102337236099 ldsub = -1.63363464867908e-07 wdsub = -1.09483094466796e-06 pdsub = 2.51546409749746e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -2.52252066206174 lpclm = 2.16706311148054e-06 wpclm = 5.18020458636356e-06 ppclm = -3.33684076576209e-12
+ pdiblc1 = 0.268689147837944 lpdiblc1 = 2.23868403869856e-07 wpdiblc1 = 1.86793964915725e-07 ppdiblc1 = -3.44711672805188e-13
+ pdiblc2 = 0.00260445737398027 lpdiblc2 = -2.46408179326341e-09 wpdiblc2 = -2.02399620662533e-09 ppdiblc2 = 3.79418328893983e-15
+ pdiblcb = -0.025
+ drout = 1.05620020214218 ldrout = -1.23425300839387e-06 wdrout = -7.6404708645772e-07 pdrout = 1.90049784531284e-12
+ pscbe1 = 29912953.3417089 lpscbe1 = -3.86788832667526 wpscbe1 = 290.10033288725 ppscbe1 = 5.95575897386117e-6
+ pscbe2 = 1.48012585562893e-08 lpscbe2 = 1.19168315419158e-15 wpscbe2 = 2.83175326807935e-16 ppscbe2 = -1.83494895409158e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -0.00104951026033924 lalpha0 = 8.37160661704906e-10 walpha0 = 1.64705990213551e-09 palpha0 = -1.28905663825057e-15
+ alpha1 = 0.0
+ beta0 = -9.50864511392075 lbeta0 = 1.83835965966143e-05 wbeta0 = 7.23363811440187e-05 pbeta0 = -2.83069885050804e-11
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -6.9913404370363e-08 lagidl = 9.05836045686824e-14 wagidl = 1.48952603932347e-13 pagidl = -1.59171639389924e-19
+ bgidl = 1524633757.17232 lbgidl = 124.06890362141 wbgidl = 141.117164835412 pbgidl = -0.000235725058334463
+ cgidl = 2756.63971351018 lcgidl = -0.00151465166819418 wcgidl = -0.00155656332138572 pcgidl = 7.56945187319887e-10
+ egidl = -2.75165686252966 legidl = 4.62699043452344e-06 wegidl = 5.61034516905343e-06 pegidl = -7.12462136311746e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.552908745121599 lkt1 = 2.79288126849516e-08 wkt1 = -4.36459100807411e-08 pkt1 = -6.82500168897112e-14
+ kt2 = -0.019032
+ at = 1644827.12968117 lat = -1.46619603088315 wat = -1.70475007975414 pat = 1.54698638282999e-6
+ ute = -1.557117677608 lute = 2.52771299464757e-07 wute = 2.01251764659688e-07 pute = -3.41250084448554e-13
+ ua1 = -3.08991162940673e-10 lua1 = 7.53372711107913e-16 wua1 = 1.3263666671314e-15 pua1 = -1.16004028707312e-21
+ ub1 = -1.04923665929664e-17 lub1 = 6.03602268220842e-24 wub1 = 8.7159866069641e-24 pub1 = -7.6230018864508e-30
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.81e-6
+ sbref = 2.81e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.61 pmos
* DC IV MOS Parameters
+ lmin = 8.0e-07 lmax = 1e-06 wmin = 1e-06 wmax = 1.5e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.40028558791717+0*(0.0/sqrt(l*w*mult))} lvth0 = 3.76537831008922e-07 wvth0 = 5.15282054326991e-07 pvth0 = -3.47609273848989e-13
+ k1 = 0.461012839457921 lk1 = 7.82179545016875e-08 wk1 = 2.08364502646493e-07 pk1 = -1.40562693485324e-13
+ k2 = -0.0396221996882736 lk2 = 5.01050647937093e-08 wk2 = 3.07687156053178e-08 pk2 = -2.07565755473474e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1426811.87145794 lvsat = -0.926426002025524 wvsat = -1.46255637388546 pvsat = 9.86640529823129e-7
+ ua = 2.2952414084009e-08 lua = -1.45579397666525e-14 wua = -2.44237861505339e-14 pua = 1.64762861371502e-20
+ ub = -1.39138910868883e-17 lub = 9.79219750921486e-24 wub = 1.72169572106126e-23 pub = -1.16145593342793e-29
+ uc = 6.87587289055318e-12 luc = -5.91339329274718e-18 wuc = -1.06242833423914e-17 puc = 7.16714154277726e-24
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0753756165271424 lu0 = -4.08251841092103e-08 wu0 = -6.47834364948746e-08 pu0 = 4.37029062594424e-14
+ a0 = 1.50385850364907 la0 = -4.77514600561664e-07 wa0 = -4.94893699766957e-07 pa0 = 3.33855289862791e-13
+ keta = 0.883520313327153 lketa = -6.39613431570498e-07 wketa = -1.08961892162516e-06 pketa = 7.35056924528331e-13
+ a1 = 0.0
+ a2 = 0.5
+ ags = -7.5765708377533 lags = 5.60748226020838e-06 wags = 8.28592741458147e-06 pags = -5.58968663387667e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.327101815135998+0*(0.009/sqrt(l*w*mult))} lvoff = 1.64256150173544e-07 wvoff = 2.71230173543555e-07 pvoff = -1.82971875072482e-13
+ nfactor = {-1.36448073131024+0*(0.02/sqrt(l*w*mult))} lnfactor = 2.16374626334189e-06 wnfactor = 3.23665128640527e-06 pnfactor = -2.18344495780899e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -1.1865e-05 lcit = 1.4750129e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.694749283603729 leta0 = -4.64074261399075e-07 weta0 = -5.6653300054246e-07 peta0 = 3.82183162165944e-13
+ etab = -0.921733775699694 letab = 6.19039455387013e-07 wetab = 9.69200762624591e-07 petab = -6.5382283446655e-13
+ dsub = 3.84682865213506 ldsub = -2.41616276255831e-06 wdsub = -3.52996367228426e-06 pdsub = 2.38131349332297e-12
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -4.08366031079326 lpclm = 3.53243584826114e-06 wpclm = 5.9688308273574e-06 ppclm = -4.0265732761353e-12
+ pdiblc1 = 0.762525815764607 lpdiblc1 = -2.08041145898804e-07 wpdiblc1 = -9.06708355449476e-07 ppdiblc1 = 6.11665456586216e-13
+ pdiblc2 = -0.0232049925472013 lpdiblc2 = 2.0108863107802e-08 wpdiblc2 = 1.01199810331266e-08 ppdiblc2 = -6.82693920494721e-15
+ pdiblcb = -0.025
+ drout = -3.39449139374158 ldrout = 2.65832186136607e-06 wdrout = 6.1613113174846e-06 pdrout = -4.15642061477512e-12
+ pscbe1 = -1132897054.29008 lpscbe1 = 1013.12574434809 wpscbe1 = 1298.38755058525 ppscbe1 = -0.00087589224162481
+ pscbe2 = 2.5201576530611e-08 lpscbe2 = -7.90443494615022e-15 wpscbe2 = -7.93641906632678e-15 ppscbe2 = 5.35390830214403e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -0.000513178058459968 lalpha0 = 3.68084517941294e-10 walpha0 = 7.57309760785761e-10 palpha0 = -5.10881164626074e-16
+ alpha1 = 0.0
+ beta0 = -109.704090392104 lbeta0 = 0.000106014533036913 wbeta0 = 0.000174792052217392 pbeta0 = -1.17914718425853e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.21028415931814e-07 lagidl = -7.6414111467602e-14 wagidl = -1.44488459953466e-13 pagidl = 9.7471915084608e-20
+ bgidl = 1254620138.2216 lbgidl = 360.222814755709 wbgidl = -561.519929847069 pbgidl = 0.00037880134467483
+ cgidl = 2761.29712620912 lcgidl = -0.00151872504134067 wcgidl = -0.0030221254678203 pcgidl = 2.03872584059157e-9
+ egidl = 10.555137049945 legidl = -7.01113152132691e-06 wegidl = -1.10890673913166e-05 pegidl = 7.48068486218219e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.117819378992 lkt1 = -3.52600346931997e-07 wkt1 = -5.32113649231635e-07 pkt1 = 3.58963867771661e-13
+ kt2 = -0.019032
+ at = -205611.11632 lat = 0.152197259069472 wat = 0.280059815385071 pat = -1.88928351458769e-7
+ ute = -0.554053706856003 lute = -6.24508449354942e-07 wute = -8.26176455385956e-07 pute = 5.57338636803367e-13
+ ua1 = 5.524e-10
+ ub1 = -3.5909e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.41e-6
+ sbref = 2.41e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.62 pmos
* DC IV MOS Parameters
+ lmin = 6e-07 lmax = 8.0e-07 wmin = 1e-06 wmax = 1.5e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.834553503+0*(0.0/sqrt(l*w*mult))} lvth0 = -5.10503347620034e-9
+ k1 = 0.45738453 lk1 = 8.0665612062e-8
+ k2 = 0.046274496373 lk2 = -7.84084636922579e-9
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 26482.8332000001 lvsat = 0.01823596718328
+ ua = 1.77765935979e-09 lua = -2.73450229694334e-16
+ ub = 5.8565225e-19 lub = 1.08055741499998e-26
+ uc = 1.604763834e-13 luc = -1.38318680902164e-18
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0177165158 lu0 = -1.92835475867999e-9
+ a0 = 0.686852 la0 = 7.36379867999997e-8
+ keta = -0.095781609 lketa = 2.10236452314e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.767854702459999 lags = -2.16672092195163e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.092270393049+0*(0.009/sqrt(l*w*mult))} lvoff = 5.83887283365537e-9
+ nfactor = {1.70823106+0*(0.02/sqrt(l*w*mult))} lnfactor = 9.08948889239981e-8
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -0.019406467399999 leta0 = 1.769520822804e-8
+ etab = -0.0138107485 letab = 6.5545812381e-9
+ dsub = 0.24951165228 ldsub = 1.05872855439121e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.2779958078 lpclm = -8.45373693418804e-8
+ pdiblc1 = 0.5860217405 lpdiblc1 = -8.89714967252998e-8
+ pdiblc2 = 0.0036505636091 lpdiblc2 = 1.99210492476115e-9
+ pdiblcb = -0.025
+ drout = 0.31784347291 ldrout = 1.53980760322914e-7
+ pscbe1 = 441057787.39 lpscbe1 = -48.6641918492942
+ pscbe2 = 1.0800700078e-08 lpscbe2 = 1.81039630878118e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.9101199429e-05 lalpha0 = -4.4830694306034e-12
+ alpha1 = 0.0
+ beta0 = 45.721312944 lbeta0 = 1.16455594637762e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -8.53727104e-08 lagidl = 6.282408835584e-14 pagidl = -1.20370621524202e-35
+ bgidl = 2357645400 lbgidl = -383.878026840001
+ cgidl = -572.088 lcgidl = 0.0007299765648
+ egidl = -2.33210108957 legidl = 1.68259932758992e-06 pegidl = -1.0097419586829e-28
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.609698460000001 lkt1 = -2.0778718884e-8
+ kt2 = -0.019032
+ at = 43730.0 lat = -0.016008258
+ ute = -1.8086978 lute = 2.2187445588e-7
+ ua1 = 5.533492e-10 lua1 = -6.40330320000525e-19
+ ub1 = -7.6755449e-18 lub1 = 2.75550144954e-24
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.02e-6
+ sbref = 2.01e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.63 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 6e-07 wmin = 1e-06 wmax = 1.5e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.023/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.678764853070431+0*(0.0/sqrt(l*w*mult))} lvth0 = -7.90423267327725e-08 wvth0 = -1.01647700387569e-07 pvth0 = 4.82419986039402e-14
+ k1 = 0.522508079695841 lk1 = 4.97579753763542e-08 wk1 = 3.73411955754665e-07 pk1 = -1.77221314201164e-13
+ k2 = 0.00865929967716889 lk2 = 1.00113259826156e-08 wk2 = -8.03973093939173e-08 pk2 = 3.81565630383532e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 214606.878350348 lvsat = -0.0710477046450755 wvsat = -0.279230095433324 pvsat = 1.32522603292656e-7
+ ua = -5.02302434896099e-09 lua = 2.95415425847889e-15 wua = 6.2138929376846e-15 pua = -2.94911358822511e-21
+ ub = 8.26864351657696e-18 lub = -3.63554208096743e-24 wub = -8.66992269130601e-24 pub = 4.11474530929384e-30
+ uc = -1.7081896607563e-11 luc = 6.80004341248943e-18 wuc = 2.73448063798356e-17 puc = -1.297784510787e-23
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0076512237337856 lu0 = 2.84863285594535e-09 wu0 = 4.30869176058705e-09 pu0 = -2.04490510957461e-15
+ a0 = 0.203698498933278 la0 = 3.02942638406265e-07 wa0 = 1.13606958976949e-06 pa0 = -5.39178627304601e-13
+ keta = 0.244580633493816 lketa = -1.40512275056165e-07 wketa = -4.75317553895164e-07 pketa = 2.25585711078645e-13
+ a1 = 0.0
+ a2 = 0.5
+ ags = -5.43373733350782 lags = 2.92160837105081e-06 wags = 8.76296200460565e-06 pags = -4.15890176738584e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.203744432699743+0*(0.009/sqrt(l*w*mult))} lvoff = 5.87444520518981e-08 wvoff = 2.58076673994774e-07 pvoff = -1.2248318947792e-13
+ nfactor = {0.514223207949755+0*(0.02/sqrt(l*w*mult))} lnfactor = 6.57571015507046e-07 wnfactor = 8.01522225619232e-07 pnfactor = -3.80402448278888e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -2.895075816e-05 lcit = 1.8486029822736e-11 wcit = 5.99762216117353e-11 pcit = -2.84647147769296e-17
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.619472441380848 leta0 = -2.8551672187935e-07 weta0 = -1.16520603822847e-06 peta0 = 5.53006785743233e-13
+ etab = 0.075831357777008 letab = -3.5989562400968e-08 wetab = -3.62136426091658e-08 petab = 1.71869947823101e-14
+ dsub = 0.300635910974266 ldsub = -1.36762876323872e-08 wdsub = -5.48147879322727e-08 pdsub = 2.60150983526566e-14
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -1.72820439814211 lpclm = 1.34220524839825e-06 wpclm = 4.7288502630379e-06 ppclm = -2.24431233483779e-12
+ pdiblc1 = 0.769030162713789 lpdiblc1 = -1.75827293907965e-07 wpdiblc1 = 6.49861553554069e-07 ppdiblc1 = -3.08424293316761e-13
+ pdiblc2 = 0.00863786686825548 lpdiblc2 = -3.7486920203405e-10 wpdiblc2 = 2.16532500746933e-08 ppdiblc2 = -1.02766324854495e-14
+ pdiblcb = -1.5830303264 lpdiblcb = 7.3944119290944e-07 wpdiblcb = 2.39904886446941e-06 ppdiblcb = -1.13858859107718e-12
+ drout = -0.697707274340001 ldrout = 6.35961144967765e-7
+ pscbe1 = 3903948901.60976 lpscbe1 = -1692.15231465799 wpscbe1 = -5504.81578096127 ppscbe1 = 0.00261258556964422
+ pscbe2 = -5.65002624059313e-08 lpscbe2 = 3.37514331036551e-14 wpscbe2 = 1.08723192412584e-13 ppscbe2 = -5.16000271190126e-20
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -3.79316146256836e-05 lalpha0 = 3.20767041197495e-11 walpha0 = 1.70204495714227e-10 palpha0 = -8.07790536659719e-17
+ alpha1 = 0.0
+ beta0 = -4.88441334303616 lbeta0 = 2.5182033642205e-05 wbeta0 = 9.44569352641404e-05 pbeta0 = -4.4829261476361e-11
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 2.21922142765006e-07 lagidl = -8.30180489562721e-14 wagidl = -4.71137211248826e-14 pagidl = 2.23601720458693e-20
+ bgidl = 3828950666.2144 lbgidl = -1082.15950618535 wbgidl = -4308.69176058707 pbgidl = 0.00204490510957462
+ cgidl = 1153.6056736 lcgidl = -8.90376526905606e-05 wcgidl = 0.00239904886446942 pcgidl = -1.13858859107719e-9
+ egidl = -0.596744115477509 legidl = 8.58998907685628e-07 wegidl = 6.08079886463889e-06 pegidl = -2.88594714115762e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.494695451039998 lkt1 = -7.53591469364165e-08 wkt1 = -3.59857329670412e-07 pkt1 = 1.70788288661577e-13
+ kt2 = -0.019032
+ at = -2430.60652799997 lat = 0.00589956585818879 wat = 0.0479809772893883 pat = -2.27717718215437e-8
+ ute = -0.883169651398397 lute = -2.1738120344632e-07 wute = -9.4522525260095e-07 pute = 4.4860390488441e-13
+ ua1 = 5.52e-10
+ ub1 = -7.81761599999998e-19 lub1 = -5.1628810464e-25
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 1.81e-6
+ sbref = 1.81e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.64 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 7.5e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.967419564992+0*(0.0/sqrt(l*w*mult))} wvth0 = 5.8431923696422e-8
+ k1 = 0.62854151472 wk1 = -4.54302622397975e-8
+ k2 = 0.00909036325278399 wk2 = 1.52776059080042e-8
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -236375.281696 wvsat = 0.329127960582374
+ ua = 1.98684992403248e-09 wua = 2.74784202053364e-16
+ ub = 5.7575184064e-19 wub = -4.4990084717011e-25
+ uc = -8.4502285941088e-11 wuc = 4.09614157831275e-17
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0157993246576 wu0 = 2.41801995912616e-9
+ a0 = 1.0066391110192 wa0 = -1.0264118604652e-7
+ keta = -0.0097115768928 wketa = 1.59055191442586e-9
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.0935404352099199 wags = 2.43727608329461e-8
+ b0 = -2.96230365312e-07 wb0 = 3.08019148929956e-13
+ b1 = -9.76977652e-10 wb1 = 1.01585745463899e-15
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.10340382694576+0*(0.009/sqrt(l*w*mult))} wvoff = -4.44648281058656e-9
+ nfactor = {1.3141095504+0*(0.02/sqrt(l*w*mult))} wnfactor = 4.16854683892282e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -1.079592e-05 wcit = 1.642453443232e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.080000000000001
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -2.7958082823 wpclm = 2.99392572832741e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0102242042336544 wpdiblc2 = -7.05619876692331e-9
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 221928871.91584 wpscbe1 = 2.89971870495731
+ pscbe2 = 1.5012430699376e-08 wpscbe2 = -1.42532109803593e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.000207239907665792 walpha0 = -1.48687985890024e-10
+ alpha1 = 0.0
+ beta0 = 43.313749698928 wbeta0 = -4.44437061545853e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -1.41191872e-08 wagidl = 3.54769943738112e-14
+ bgidl = 947008104.0 wbgidl = 596.210599893217
+ cgidl = 2031.8368 wcgidl = -0.0006569813772928
+ egidl = 2.8810904770144 wegidl = -1.41532381241846e-6
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.524408160000001 wkt1 = -3.28490688646398e-8
+ kt2 = -0.019032
+ at = -481852.5144 wat = 0.658131094703063
+ ute = -2.0163931088 wute = 4.78610933357804e-7
+ ua1 = 2.2096e-11
+ ub1 = -5.2151516496e-18 wub1 = 2.22355347144748e-24
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.65 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 7.5e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.0042960313325+0*(0.0/sqrt(l*w*mult))} lvth0 = 7.3290501793091e-07 wvth0 = 9.67759258914085e-08 pvth0 = -7.62071706024482e-13
+ k1 = 0.657212614871176 lk1 = -5.69826647064562e-07 wk1 = -7.52423574925894e-08 pk1 = 5.92503468311143e-13
+ k2 = -0.000551354568401607 lk2 = 1.91625285008935e-07 wk2 = 2.53030255316017e-08 pk2 = -1.99251204851151e-13
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -444088.384266277 lvsat = 4.12821482834323 wvsat = 0.545107213782538 pvsat = -4.29250126565197e-6
+ ua = 1.81343324121766e-09 lua = 3.44658720427142e-15 wua = 4.55102175177481e-16 pua = -3.58374758865259e-21
+ ub = 8.59684875831979e-19 lub = -5.6430555012265e-24 wub = -7.45133281430588e-25 pub = 5.86762653795331e-30
+ uc = -1.10353091028962e-10 luc = 5.13774410799467e-16 wuc = 6.78409795102789e-17 puc = -5.34220577251643e-22
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0142733089799948 lu0 = 3.03289511861334e-08 wu0 = 4.00476495663738e-09 pu0 = -3.15359221275367e-14
+ a0 = 1.07141610282352 la0 = -1.28741680131406e-06 wa0 = -1.69996043016681e-07 pa0 = 1.33865084033915e-12
+ keta = -0.0107153763644703 lketa = 1.99501129796574e-08 wketa = 2.63429858987071e-09 pketa = -2.07440476757958e-14
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.0781587527729229 lags = 3.05704785762341e-07 wags = 4.03665727042058e-08 pags = -3.1787061341654e-13
+ b0 = -4.90621668202489e-07 lb0 = 3.86344938842733e-12 wb0 = 5.10146448110276e-13 pb0 = -4.01719922028918e-18
+ b1 = -1.61808667020327e-09 lb1 = 1.27417852931826e-14 wb1 = 1.68248004733068e-15 pb1 = -1.32488573807101e-20
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.10059764560985+0*(0.009/sqrt(l*w*mult))} lvoff = -5.57717315786739e-08 wvoff = -7.3643389389403e-09 pvoff = 5.79912234085794e-14
+ nfactor = {1.05103199369832+0*(0.02/sqrt(l*w*mult))} lnfactor = 5.22856120842322e-06 wnfactor = 6.90401675040462e-07 pnfactor = -5.43663703027362e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -2.11614659693333e-05 lcit = 2.06011079922112e-10 wcit = 2.72025876690489e-11 pcit = -2.14209496858693e-16
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.080000000000001
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -4.68527887238746 lpclm = 3.75524721897523e-05 wpclm = 4.958589690018e-06 ppclm = -3.90469103730157e-11
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0146773808511523 lpdiblc2 = -8.8505104002124e-08 wpdiblc2 = -1.16865940010912e-08 ppdiblc2 = 9.20272531209926e-14
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 220098855.506046 lpscbe1 = 36.3708441380895 wpscbe1 = 4.80256244779525 ppscbe1 = -3.78182582514083e-5
+ pscbe2 = 1.50214259201682e-08 lpscbe2 = -1.78776415156389e-16 wpscbe2 = -2.36064055792064e-17 ppscbe2 = 1.85891001373978e-22
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.000301077097339662 lalpha0 = -1.86497660989231e-09 walpha0 = -2.46259520364156e-10 palpha0 = 1.93919521905958e-15
+ alpha1 = 0.0
+ beta0 = 46.1185980256262 lbeta0 = -5.57452385537959e-05 wbeta0 = -7.36084068616601e-06 pbeta0 = 5.7963676067283e-11
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -3.650876649376e-08 lagidl = 4.44983932631763e-13 wagidl = 5.87575893651457e-14 pagidl = -4.62692513214776e-19
+ bgidl = 570738785.3132 lbgidl = 7478.20220117268 wbgidl = 987.453932386476 pbgidl = -0.00777580473597055
+ cgidl = 2446.45863877333 lcgidl = -0.00824044319688449 wcgidl = -0.00108810350676196 pcgidl = 8.56837987434771e-9
+ egidl = 3.77430325571253 legidl = -1.77522466915139e-05 wegidl = -2.34408288685767e-06 pegidl = 1.84587151008494e-11
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.503677068061334 lkt1 = -4.1202215984422e-07 wkt1 = -5.44051753380975e-08 pkt1 = 4.28418993717383e-13
+ kt2 = -0.019032
+ at = -897199.941391186 lat = 8.25486397247904 wat = 1.09000768789879 pat = -8.58337453912782e-6
+ ute = -2.31844511834637 lute = 6.00316286893035e-06 wute = 7.92683404676086e-07 pute = -6.24206473846231e-12
+ ua1 = 2.2096e-11
+ ub1 = -6.61843926292834e-18 lub1 = 2.78897799998556e-23 wub1 = 3.68268631863584e-24 pub1 = -2.89996816847298e-29
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.66 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 7.5e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.925593902757065+0*(0.0/sqrt(l*w*mult))} lvth0 = 1.13157236250774e-07 wvth0 = -2.25916678945701e-09 pvth0 = 1.77900348002583e-14
+ k1 = 0.460945144239072 lk1 = 9.75701177175007e-07 wk1 = 1.0844000589394e-07 pk1 = -8.53921670412419e-13
+ k2 = 0.0620520405221855 lk2 = -3.01351409971402e-07 wk2 = -3.37826033185492e-08 pk2 = 2.66024488092247e-13
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 225314.152025792 lvsat = -1.1430623839423 wvsat = -0.19129733434107 pvsat = 1.50638998900219e-6
+ ua = 3.6514099453057e-09 lua = -1.10267441497402e-14 wua = -1.16994115661925e-15 pua = 9.21281863191397e-21
+ ub = -8.05148726007466e-19 lub = 7.46684317981839e-24 wub = 8.53678673159776e-25 pub = -6.72237807966397e-30
+ uc = -6.82138008519372e-11 luc = 1.81944356371464e-16 wuc = 8.70873159775082e-18 puc = -6.85777778396487e-23
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0232192826828764 lu0 = -4.01170133345785e-08 wu0 = -4.58674496760899e-09 pu0 = 3.61187819219338e-14
+ a0 = 0.962353300724496 la0 = -4.28590859905125e-07 wa0 = -1.90816863657677e-08 pa0 = 1.50260647455875e-13
+ keta = -7.16043979827885e-05 lketa = -6.38653337476448e-08 wketa = -6.77590940584347e-09 pketa = 5.33575762072549e-14
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.162668500977929 lags = -3.59775677452798e-07 wags = -4.17605708261119e-08 pags = 3.28847791027301e-13
+ b0 = 2.86943543359469e-07 lb0 = -2.25956562653848e-12 wb0 = -2.98362748611003e-13 pb0 = 2.3494873002122e-18
+ b1 = 9.46349402609802e-10 lb1 = -7.45212300579114e-15 wb1 = -9.84010323436061e-16 pb1 = 7.7486876929296e-21
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.154566456747719+0*(0.009/sqrt(l*w*mult))} lvoff = 3.69211068607584e-07 wvoff = 3.80661935584135e-08 pvoff = -2.99756047795083e-13
+ nfactor = {1.87156572575559+0*(0.02/sqrt(l*w*mult))} lnfactor = -1.23281371803499e-06 wnfactor = -2.20730141105123e-07 pnfactor = 1.73816156914641e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.56749999999995e-07 lcit = 3.813865645e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.080000000000001
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.47166228843676 lpclm = 4.37192703777412e-06 wpclm = -2.587784236074e-07 ppclm = 2.03777657453883e-12
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00551879131209 lpdiblc2 = -1.63848748178239e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 226044860.806281 lpscbe1 = -10.451569199141 wpscbe1 = -1.72358516410304 ppscbe1 = 1.3572543733245e-5
+ pscbe2 = 1.49505315118213e-08 lpscbe2 = 3.79488692812166e-16 wpscbe2 = 4.13809353477399e-17 ppscbe2 = -3.2585831348931e-22
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.000184548275490656 lalpha0 = -9.47358749360117e-10 walpha0 = -6.03883333092269e-11 palpha0 = 4.75533969476838e-16
+ alpha1 = -4.02879358160001e-10 lalpha1 = 3.17251379376674e-15 walpha1 = 3.18192505557336e-16 palpha1 = -2.5056387042618e-21
+ beta0 = 180.094822369448 lbeta0 = -0.00111075441477166 wbeta0 = -0.000110369878441321 pbeta0 = 8.69118644774025e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -1.74204202848001e-09 lagidl = 1.71209884157469e-13 wagidl = 8.90939015560543e-15 pagidl = -7.01578837193304e-20
+ bgidl = 2269601031.33536 lbgidl = -5899.65844135344 wbgidl = -730.569992759642 pbgidl = 0.00575294646498508
+ cgidl = 4446.1158557728 lcgidl = -0.0239869439178685 wcgidl = -0.00225280293934594 pcgidl = 1.77399220261735e-8
+ egidl = -1.73262984407209 legidl = 2.56126486960501e-05 wegidl = 2.89848362631796e-06 pegidl = -2.28243991638034e-11
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.506025564184 lkt1 = -3.93528692276676e-07 wkt1 = -3.18192505557337e-08 pkt1 = 2.5056387042618e-13
+ kt2 = -0.019032
+ at = 487975.678619065 lat = -2.65283996485369 wat = -0.419345903074013 pat = 3.30218124834662e-6
+ ute = -1.697232305 lute = 1.111360448953e-6
+ ua1 = 2.2096e-11
+ ub1 = -3.732379185e-18 lub1 = 5.16321131020101e-24
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.67 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 7.5e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.861626567137496+0*(0.0/sqrt(l*w*mult))} lvth0 = -1.346906023408e-07 wvth0 = -4.79930431180489e-08 pvth0 = 1.94990512023022e-13
+ k1 = 0.724959302111809 lk1 = -4.72480789186998e-08 wk1 = -1.13304361709554e-07 pk1 = 5.24905630407679e-15
+ k2 = -0.0209702915102319 lk2 = 2.03269177214029e-08 wk2 = 3.39387714452409e-08 pk2 = 3.63124943246637e-15
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -104039.705453315 lvsat = 0.133052072246247 wvsat = 0.329840055470427 pvsat = -5.12808941561435e-7
+ ua = 1.13762628426069e-09 lua = -1.28683797665525e-15 wua = 1.16975143172155e-15 pua = 1.47445729128688e-22
+ ub = -5.36788081746109e-19 lub = 6.42705302756334e-24 wub = 6.58656574687875e-25 pub = -5.96674545692474e-30
+ uc = -1.44190891242425e-12 luc = -7.67700161373727e-17 wuc = -4.67306453106914e-17 puc = 1.46227631929802e-22
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.00999305325479524 lu0 = 1.11293352074649e-08 wu0 = 8.55000393221974e-09 pu0 = -1.47808653653426e-14
+ a0 = 0.186974286263501 la0 = 2.57569266952546e-06 wa0 = 6.46396290994706e-07 pa0 = -2.42820032362501e-12
+ keta = 0.305656703778136 lketa = -1.24844023660684e-06 wketa = -2.25654359257137e-07 pketa = 9.01424018001078e-13
+ a1 = 0.0
+ a2 = 0.5
+ ags = -1.2509419261581 lags = 5.11739928352846e-06 wags = 8.58218418514019e-07 pags = -3.15821080106997e-12
+ b0 = -1.2575373400025e-07 lb0 = -6.60528755680508e-13 wb0 = 1.30758229598524e-13 pb0 = 6.8681515804157e-19
+ b1 = -8.5512825683432e-10 lb1 = -4.72117666508944e-16 wb1 = 8.89158940943299e-16 pb1 = 4.90906061165333e-22
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.00321545258693534+0*(0.009/sqrt(l*w*mult))} lvoff = -2.17213532113787e-07 wvoff = -1.0822576413508e-07 pvoff = 2.67066771484127e-13
+ nfactor = {1.8580001097103+0*(0.02/sqrt(l*w*mult))} lnfactor = -1.18025238210591e-06 wnfactor = -1.330397340833e-07 pnfactor = 1.39839631809964e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 2.19058027878373e-05 lcit = -4.61302234817545e-11 wcit = -9.40315541862276e-12 pcit = 3.64334659849958e-17
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.332650189792001 leta0 = -9.78918425368083e-07 weta0 = -1.84736593480962e-07 peta0 = 7.15780405101337e-13
+ etab = -0.133084834750246 letab = 2.44428500723305e-07 wetab = -1.99515520959438e-09 petab = 7.73042837509446e-15
+ dsub = 1.0068806298801 ldsub = -1.73148368853344e-06 wdsub = -1.7228445418681e-07 pdsub = 6.67533346192216e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -2.68179337095536 lpclm = 1.29353009301007e-05 wpclm = 2.77372946868167e-06 ppclm = -9.7119785049244e-12
+ pdiblc1 = 0.850226524828679 lpdiblc1 = -1.7831936931012e-06 wpdiblc1 = -4.79426929509046e-07 ppdiblc1 = 1.85758758107575e-12
+ pdiblc2 = 0.00348315467889863 lpdiblc2 = -8.49759711886063e-09 wpdiblc2 = -2.28043346250008e-09 ppdiblc2 = 8.83576749380281e-15
+ pdiblcb = -0.025
+ drout = -0.141333179345208 ldrout = 2.71738553669095e-06 wdrout = 6.53224407185896e-07 pdrout = -2.53098328808248e-12
+ pscbe1 = 48157133.9314482 lpscbe1 = 678.792217350087 wpscbe1 = 101.252665277451 ppscbe1 = -0.0003854192362276
+ pscbe2 = 1.45594916822818e-08 lpscbe2 = 1.89461161634587e-15 wpscbe2 = 6.99117287553356e-16 ppscbe2 = -2.87432358374517e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -0.0013627359091259 lalpha0 = 5.0477485523552e-09 walpha0 = 1.1053219976391e-09 palpha0 = -4.04112727881556e-15
+ alpha1 = 1.10186903264e-09 lalpha1 = -2.65778432122694e-15 walpha1 = -9.44279333582941e-16 palpha1 = 2.38593468367112e-21
+ beta0 = -413.347629918581 lbeta0 = 0.00118859771086354 wbeta0 = 0.00038190254472155 pbeta0 = -1.03824008601283e-9
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -7.33933499770058e-08 lagidl = 4.48830041934828e-13 wagidl = 1.05013812271571e-13 pagidl = -4.42524077649851e-19
+ bgidl = -1766712658.15343 lbgidl = 9739.44257993987 wbgidl = 3237.99812048367 pbgidl = -0.00962366754658748
+ cgidl = -1709.6280860896 lcgidl = -0.000135898440728436 wcgidl = 0.00195008300220522 pcgidl = 1.45542015703939e-9
+ egidl = 6.46309143128607 legidl = -6.14249295745266e-06 wegidl = -4.1115650003768e-06 pegidl = 4.33673524518813e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.6983645760176 lkt1 = 3.51708042973794e-07 wkt1 = 1.65243627525996e-07 pkt1 = -5.12975956989291e-13
+ kt2 = -0.019032
+ at = -343651.825814402 lat = 0.56938396382423 wat = 0.783381670059825 pat = -1.35790700651775e-6
+ ute = -1.5527969255072 lute = 5.51731127570197e-07 wute = 1.41631388335406e-07 pute = -5.4876497724436e-13
+ ua1 = -1.33634910214067e-09 lua1 = 5.26343139275424e-15 wua1 = 6.80323294925891e-16 pua1 = -2.63598063851986e-21
+ ub1 = -4.363120468928e-18 lub1 = 7.60708148890843e-24 wub1 = 2.43236514749934e-24 pub1 = -9.42444200050093e-30
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.68 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 7.5e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.941633344352694+0*(0.0/sqrt(l*w*mult))} lvth0 = 1.52901022268087e-08 wvth0 = 4.34433094426981e-08 pvth0 = 2.3583925512644e-14
+ k1 = 0.689605983469344 lk1 = 1.90252522084631e-08 wk1 = -1.02488654680154e-07 pk1 = -1.50260680932357e-14
+ k2 = -0.0130560132643047 lk2 = 5.49081172158777e-09 wk2 = 3.8868843591055e-08 pk2 = -5.61066381207687e-15
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -36854.758557664 lvsat = 0.00710717079565937 wvsat = 0.037637957229444 pvsat = 3.49531118011113e-8
+ ua = 3.05508005493699e-09 lua = -4.88129681516504e-15 wua = -8.079929974722e-16 pua = 3.8549254360953e-21
+ ub = 7.59977443032097e-19 lub = 3.99613637481411e-24 wub = -8.57642522668523e-25 pub = -3.12429116902044e-30
+ uc = -7.91187129994723e-11 luc = 6.88429208042077e-17 wuc = 6.02785808758452e-17 puc = -5.437186347948e-23
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0225524397886685 lu0 = -1.24144907889339e-08 wu0 = -4.29270718718999e-09 pu0 = 9.29408089910287e-15
+ a0 = 1.88052437097126 la0 = -5.99036319267711e-07 wa0 = -9.01302851455618e-07 pa0 = 4.73116488812361e-13
+ keta = -0.447539623549705 lketa = 1.63501598601936e-07 wketa = 3.20938600335896e-07 pketa = -1.23219144052022e-13
+ a1 = 0.0
+ a2 = 0.5
+ ags = 1.57658563834099 lags = -1.8308388888153e-07 wags = -9.0365596758064e-07 pags = 1.44598923103077e-13
+ b0 = -2.3883317309376e-07 lb0 = -4.48550039155813e-13 wb0 = 2.483377780502e-13 pb0 = 4.66400536514058e-19
+ b1 = -1.28298259579168e-09 lb1 = 3.29938077300523e-16 wb1 = 1.33404017117381e-15 pb1 = -3.43068293024775e-22
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.142779103231042+0*(0.009/sqrt(l*w*mult))} lvoff = 4.44124873836564e-08 wvoff = 5.29518611555364e-08 pvoff = -3.50768048856624e-14
+ nfactor = {1.1214632177441+0*(0.02/sqrt(l*w*mult))} lnfactor = 2.0045967557394e-07 wnfactor = 7.20983537306038e-07 pnfactor = -2.02555706446808e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 4.37650605632534e-06 lcit = -1.32698038288621e-11 wcit = 4.44141302273848e-12 pcit = 1.048043798482e-17
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -0.399395742385877 leta0 = 3.93374879092568e-07 weta0 = 3.79330379842239e-07 peta0 = -3.41619543090337e-13
+ etab = -0.014186028343589 letab = 2.15407982333848e-08 wetab = 1.42024311947044e-08 petab = -2.2633567098404e-14
+ dsub = -0.0910659284626156 ldsub = 3.26726929735816e-07 wdsub = 3.2146406197122e-07 pdsub = -2.58047622197628e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 6.53054514013444 lpclm = -4.33414884278825e-06 wpclm = -4.23313702249682e-06 ppclm = 3.42309341943879e-12
+ pdiblc1 = 0.137830874897232 lpdiblc1 = -4.47736807739711e-07 wpdiblc1 = 3.22859873686386e-07 ppdiblc1 = 3.53620739805593e-13
+ pdiblc2 = -0.00367877890980694 lpdiblc2 = 4.92816358652682e-09 wpdiblc2 = 4.50928774831148e-09 ppdiblc2 = -3.89224388798454e-15
+ pdiblcb = -0.025
+ drout = -0.0085691123958771 ldrout = 2.46850601678773e-06 wdrout = 3.43095787721693e-07 pdrout = -1.94961617803488e-12
+ pscbe1 = 406130269.905382 lpscbe1 = 7.73577665335051 wpscbe1 = -101.088928006391 ppscbe1 = -6.10968545770949e-6
+ pscbe2 = 1.68415667514854e-08 lpscbe2 = -2.38336630838316e-15 wpscbe2 = -1.83832897332414e-15 ppscbe2 = 1.88237317689578e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.00222313300998485 lalpha0 = -1.67432132340981e-09 walpha0 = -1.75582147977439e-09 palpha0 = 1.32237228394377e-15
+ alpha1 = -3.159184e-10 walpha1 = 3.284906886464e-16
+ beta0 = 240.319767956577 lbeta0 = -3.67671931932286e-05 wbeta0 = -0.000187434203453033 pbeta0 = 2.90385821152392e-11
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 3.04694093056246e-07 lagidl = -2.59932678775306e-13 wagidl = -2.40562773461851e-13 pagidl = 2.05293789966022e-19
+ bgidl = 3656480244.03264 lbgidl = -426.874834498147 wbgidl = -2075.568284816 pbgidl = 0.000337144036787298
+ cgidl = -1904.35608665357 lcgidl = 0.000229138669128778 wcgidl = 0.00328992146764135 pcgidl = -1.05624103026717e-9
+ egidl = 8.12290574452314 legidl = -9.25398086904687e-06 wegidl = -5.69698153150963e-06 pegidl = 7.30875707444974e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.4270816144928 lkt1 = -1.56838996700597e-07 wkt1 = -1.74480457200045e-07 pkt1 = 1.23870812238145e-13
+ kt2 = -0.019032
+ at = -101063.74884745 lat = 0.114628354741979 wat = 0.1106202721764 pat = -9.67484900454797e-8
+ ute = -1.0911469089856 lute = -3.13677993401195e-07 wute = -2.83262776670809e-07 pute = 2.4774162447629e-13
+ ua1 = 2.27518232588134e-09 lua1 = -1.50674542221582e-15 wua1 = -1.36064658985178e-15 pua1 = 1.19002150748437e-21
+ ub1 = 2.568576997856e-18 lub1 = -5.38707858232486e-24 wub1 = -4.86473029499868e-24 pub1 = 4.25469311600584e-30
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.81e-6
+ sbref = 2.81e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.69 pmos
* DC IV MOS Parameters
+ lmin = 8.0e-07 lmax = 1e-06 wmin = 7.5e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.12794076978978+0*(0.0/sqrt(l*w*mult))} lvth0 = 1.78234576514079e-07 wvth0 = 2.32099001817402e-07 pvth0 = -1.4141434303827e-13
+ k1 = 0.982257665693918 lk1 = -2.36927909065149e-07 wk1 = -3.33623782694394e-07 pk1 = 1.87124714868019e-13
+ k2 = -0.11296823545104 lk2 = 9.28740412461063e-08 wk2 = 1.07033630207299e-07 pk2 = -6.52275861866438e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -190627.247556251 lvsat = 0.141596589673823 wvsat = 0.219250352309021 pvsat = -1.23885088935486e-7
+ ua = -8.64204881923415e-09 lua = 5.34901209818504e-15 wua = 8.42800999840679e-15 pua = -4.22288278410046e-21
+ ub = 1.02876230189237e-17 lub = -4.33674244586066e-24 wub = -7.94768035055428e-24 pub = 3.07665591524844e-30
+ uc = -5.06286415199914e-12 luc = 4.07367540220764e-18 wuc = 1.78956767950632e-18 puc = -3.21737253796199e-24
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = -0.00235343610166877 lu0 = 9.36818826475503e-09 wu0 = 1.60389215123528e-08 pu0 = -8.48796156151726e-15
+ a0 = 1.93953832901333 la0 = -6.50649926971301e-07 wa0 = -9.47911839461411e-07 pa0 = 5.13880709722226e-13
+ keta = -0.580693235187344 lketa = 2.79957747340214e-07 wketa = 4.32864469266023e-07 pketa = -2.21109509018312e-13
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.265257202121692 lags = 9.63803961435867e-07 wags = 1.32025986031618e-07 pags = -7.61208513526202e-13
+ b0 = -3.28716766171808e-06 lb0 = 2.21752330459501e-12 wb0 = 3.41798378598381e-12 pb0 = -2.30577186202468e-18
+ b1 = -3.9607925048944e-09 lb1 = 2.67195062380176e-15 wb1 = 4.11841620341918e-15 pb1 = -2.77828357082657e-21
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0362979278706692+0*(0.009/sqrt(l*w*mult))} lvoff = -4.87159485865259e-08 wvoff = -3.11465452193851e-08 pvoff = 3.84756613298439e-14
+ nfactor = {1.22084322340144+0*(0.02/sqrt(l*w*mult))} lnfactor = 1.13541922626027e-07 wnfactor = 5.48441779591874e-07 pnfactor = -5.16506851499969e-14
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -8.09405581599999e-05 lcit = 6.13485005347359e-11 wcit = 7.18244890725353e-11 pcit = -4.84528003283323e-17
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.50937680878225 leta0 = -4.01437594159077e-07 weta0 = -3.73783442712985e-07 peta0 = 3.17053806116462e-13
+ etab = 0.0568557483374108 letab = -4.05923396518177e-08 wetab = -4.83327101110937e-08 petab = 3.2059667487647e-14
+ dsub = 0.88165126782402 ldsub = -5.24011530136476e-07 wdsub = -4.4678408878718e-07 pdsub = 4.13862210455668e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 3.19198305534001 lpclm = -1.41424244342705e-06 wpclm = -1.59635404217452e-06 ppclm = 1.11696302484891e-12
+ pdiblc1 = -2.18222083870968 lpdiblc1 = 1.58138042098089e-06 wpdiblc1 = 2.15522743688627e-06 ppdiblc1 = -1.24896793096902e-12
+ pdiblc2 = -0.0624491211117789 lpdiblc2 = 5.63287048763716e-08 wpdiblc2 = 5.09258689380602e-08 ppdiblc2 = -4.44881857965387e-14
+ pdiblcb = -0.025
+ drout = 9.1816192288392 ldrout = -5.56923270645647e-06 wdrout = -6.9152782034324e-06 pdrout = 4.39855771462849e-12
+ pscbe1 = -397061638.084644 lpscbe1 = 710.207419381427 wpscbe1 = 533.268828156499 ppscbe1 = -0.000560918978997774
+ pscbe2 = 2.7220025292658e-08 lpscbe2 = -1.14603661484927e-14 wpscbe2 = -1.00351940153081e-14 ppscbe2 = 9.05135134261495e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.000894836757326878 lalpha0 = -5.12593420835151e-10 walpha0 = -7.0673841261014e-10 palpha0 = 4.04844233401919e-16
+ alpha1 = -3.159184e-10 walpha1 = 3.284906886464e-16
+ beta0 = 233.411159376176 lbeta0 = -3.07249241288097e-05 wbeta0 = -0.000181977812030666 pbeta0 = 2.42664221772374e-11
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -7.34758418815743e-08 lagidl = 7.08147463213113e-14 wagidl = 5.77562893038647e-14 pagidl = -5.56160623288729e-20
+ bgidl = -277104458.419197 lbgidl = 3013.43834626623 wbgidl = 1031.16117884164 pbgidl = -0.00238000155212768
+ cgidl = -3744.17749174624 lcgidl = 0.00183824647002283 wcgidl = 0.00374224101803121 pcgidl = -1.45183970903815e-9
+ egidl = -3.32934016489497 legidl = 7.62153403330207e-07 wegidl = 3.34795647876515e-06 pegidl = -6.01945709336584e-13
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.566007877104001 lkt1 = -3.53340874208398e-08 wkt1 = -6.60890416487684e-08 pkt1 = 2.9071680196999e-14
+ kt2 = -0.019032
+ at = -42829.2763199999 lat = 0.0636964850694718 wat = 0.110799909280431 pat = -9.69056006566646e-8
+ ute = -1.34861 lute = -8.85007740000023e-8
+ ua1 = 5.524e-10
+ ub1 = -3.5909e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.41e-6
+ sbref = 2.41e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.70 pmos
* DC IV MOS Parameters
+ lmin = 6e-07 lmax = 8.0e-07 wmin = 7.5e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.850318020711041+0*(0.0/sqrt(l*w*mult))} lvth0 = -9.04973001443431e-09 wvth0 = 1.63918824578666e-08 pvth0 = 4.10167968167032e-15
+ k1 = 0.215048516870721 lk1 = 2.80631382730979e-07 wk1 = 2.51980017107772e-07 pk1 = -2.07923608478523e-13
+ k2 = 0.101376788959421 lk2 = -5.17231122211904e-08 wk2 = -5.72951434221899e-08 pk2 = 4.56286045038093e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -128278.556720906 lvsat = 0.0995361628362995 wvsat = 0.160920274194198 pvsat = -8.45356182392271e-8
+ ua = -7.08986644949028e-09 lua = 4.30190987155582e-15 wua = 9.2204178663864e-15 pua = -4.75744113183951e-21
+ ub = 1.8679272646917e-17 lub = -9.99774928490493e-24 wub = -1.88136741142327e-23 pub = 1.04068553082259e-29
+ uc = 9.14310839168304e-12 luc = -5.50967367576036e-18 wuc = -9.34010483168467e-18 puc = 4.29070453808745e-24
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0166037957831127 lu0 = -3.42036036471851e-09 wu0 = 1.15700182267939e-09 pu0 = 1.55138146113643e-15
+ a0 = 1.05307664577104 la0 = -5.26428754560552e-08 wa0 = -3.80798921774145e-07 pa0 = 1.31306335450397e-13
+ keta = -0.599232422040336 lketa = 2.92464282791243e-07 wketa = 5.23486141596089e-07 pketa = -2.82242889172174e-13
+ a1 = 0.0
+ a2 = 0.5
+ ags = 5.73630911270508 lags = -2.72696765744369e-06 wags = -5.1661790219552e-06 pags = 2.8129605848617e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.381134486453465+0*(0.009/sqrt(l*w*mult))} lvoff = 1.83910793833428e-07 wvoff = 3.00359728865589e-07 pvoff = -1.8515847116788e-13
+ nfactor = {-4.70549690904+0*(0.02/sqrt(l*w*mult))} lnfactor = 4.11145097597102e-06 wnfactor = 6.66896868729592e-06 pnfactor = -4.18055813708715e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -2.748371816e-05 lcit = 2.5286516270736e-11 wcit = 3.89754202078954e-11 pcit = -2.62928184722462e-17
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -0.308956774158697 leta0 = 1.50610240892886e-07 weta0 = 3.01073250766467e-07 peta0 = -1.38204519304776e-13
+ etab = -0.0111872591170016 letab = 5.30947317692896e-09 wetab = -2.72789376648421e-09 petab = 1.2946583815734e-15
+ dsub = -0.151150943936232 ldsub = 1.7271684191699e-07 wdsub = 4.16607364895254e-07 pdsub = -1.68581664198501e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.98096439415947 lpclm = -5.97289254594659e-07 wpclm = -7.30943924222234e-07 ppclm = 5.33157359278299e-13
+ pdiblc1 = 1.10714734006376 lpdiblc1 = -6.37627352419668e-07 wpdiblc1 = -5.41864313924e-07 ppdiblc1 = 5.70490164127581e-13
+ pdiblc2 = 0.0276209148896758 lpdiblc2 = -4.43254141020984e-09 wpdiblc2 = -2.49242753801377e-08 ppdiblc2 = 6.68032156051749e-15
+ pdiblcb = -0.025
+ drout = 4.27443425945134 ldrout = -2.25884572610742e-06 wdrout = -4.11404727348254e-06 pdrout = 2.50884732928431e-12
+ pscbe1 = 1869334996.57374 lpscbe1 = -818.703750359118 wpscbe1 = -1485.11692900042 ppscbe1 = 0.000800684052780282
+ pscbe2 = -1.18598226243546e-09 lpscbe2 = 7.70232654817333e-15 wpscbe2 = 1.24637043508555e-14 ppscbe2 = -6.12640549519897e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.000419522949745473 lalpha0 = -1.91946726240736e-10 walpha0 = -3.95561014292068e-10 palpha0 = 1.94923960496548e-16
+ alpha1 = -1.0655927632e-09 lalpha1 = 5.0573032541472e-16 walpha1 = 1.10799909280431e-15 palpha1 = -5.25856369444924e-22
+ beta0 = 529.281628838765 lbeta0 = -0.000230319142828272 wbeta0 = -0.000502804082226113 pbeta0 = 2.40695824051086e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -1.39482994072794e-07 lagidl = 1.15343171189508e-13 wagidl = 5.62636565218361e-14 pagidl = -5.46091322541165e-20
+ bgidl = 11895841096.064 lbgidl = -5198.43072478814 wbgidl = -9917.77773198457 pbgidl = 0.00500615263711568
+ cgidl = -6974.65577245792 lcgidl = 0.00401752711819093 wcgidl = 0.00665736435953066 pcgidl = -3.41838191521367e-9
+ egidl = -12.2466741222871 legidl = 6.77778689098697e-06 wegidl = 1.03091333811272e-05 pegidl = -5.29795564767e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.160269784976 lkt1 = -3.0904500437039e-07 wkt1 = -4.67314138575255e-07 pkt1 = 2.99738130583606e-13
+ kt2 = -0.019032
+ at = 150289.27632 lat = -0.066581290541472 wat = -0.110799909280431 pat = 5.25856369444924e-8
+ ute = -1.8086978 lute = 2.21874455880003e-7
+ ua1 = 5.533492e-10 lua1 = -6.40330319998947e-19
+ ub1 = -7.6755449e-18 lub1 = 2.75550144954e-24
+ uc1 = 4.31105307045504e-10 luc1 = -3.64489960132897e-16 wuc1 = -5.61807297044687e-16 puc1 = 3.78995202586346e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.02e-6
+ sbref = 2.01e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.71 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 6e-07 wmin = 7.5e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.02/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.465711229499327+0*(0.0/sqrt(l*w*mult))} lvth0 = -1.91584113123514e-07 wvth0 = -3.2318000596231e-07 pvth0 = 1.65262497925887e-13
+ k1 = 1.40891139049952 lk1 = -2.85975937093249e-07 wk1 = -5.48266661205758e-07 pk1 = 1.71873465049079e-13
+ k2 = -0.085180584053535 lk2 = 3.68170170107584e-08 wk2 = 1.71770263497336e-08 pk2 = 1.02841127300544e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -291810.137294199 lvsat = 0.177148250976385 wvsat = 0.247340291765814 pvsat = -1.25550558578716e-7
+ ua = 1.17755398093508e-08 lua = -4.65161193889015e-15 wua = -1.12531868798714e-14 pua = 4.95933168073442e-21
+ ub = -2.74717766484442e-17 lub = 1.19055387106735e-23 wub = 2.84928232346023e-23 pub = -1.20448083335312e-29
+ uc = 2.07680906036343e-11 luc = -1.10268902335524e-17 wuc = -1.20114589224186e-17 puc = 5.55852918954976e-24
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = -0.00440838821795336 lu0 = 6.55202216218741e-09 wu0 = 1.68482280295574e-08 pu0 = -5.89567449664788e-15
+ a0 = 1.31809046519232 la0 = -1.78418434153395e-07 wa0 = -2.26707191787959e-08 pa0 = -3.86613095013561e-14
+ keta = -0.352858881886385 lketa = 1.75535400634177e-07 wketa = 1.45897664439107e-07 pketa = -1.0303939791347e-13
+ a1 = 0.0
+ a2 = 0.5
+ ags = 9.85325287705503 lags = -4.68086916800417e-06 wags = -7.13238926837676e-06 pags = 3.74612396781337e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {0.618875453277678+0*(0.009/sqrt(l*w*mult))} lvoff = -2.90693923562972e-07 wvoff = -5.97280192965004e-07 pvoff = 2.4086143573292e-13
+ nfactor = {15.2980532017581+0*(0.02/sqrt(l*w*mult))} lnfactor = -5.38223390661376e-06 wnfactor = -1.45706450666227e-05 pnfactor = 5.89976255052264e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 0.00016286895264 lcit = -6.50548612909441e-11 wcit = -1.39477146399262e-10 pcit = 5.84007696395106e-17
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -1.59036930112084 leta0 = 7.58768626189116e-07 weta0 = 1.13257856625781e-06 peta0 = -5.32836942036966e-13
+ etab = 0.118798875366557 letab = -5.6381946248968e-08 wetab = -8.08910955287085e-08 petab = 3.8390913937925e-14
+ dsub = -0.13327324930543 ldsub = 1.64232088045211e-07 wdsub = 3.96362221289916e-07 pdsub = -1.58973319043408e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 5.74353615952729 lpclm = -2.38300581443822e-06 wpclm = -3.0402356818645e-06 ppclm = 1.62914722745532e-12
+ pdiblc1 = -1.05560387297936 lpdiblc1 = 3.88814373290598e-07 wpdiblc1 = 2.54710872533167e-06 ppdiblc1 = -8.95536440303157e-13
+ pdiblc2 = 0.0982357380203156 lpdiblc2 = -3.79463364680114e-08 wpdiblc2 = -7.15102579577341e-08 ppdiblc2 = 2.87900288918448e-14
+ pdiblcb = 3.09106065280001 lpdiblcb = -1.47888238581888e-06 wpdiblcb = -2.46105223933884e-06 ppdiblcb = 1.16801539279021e-12
+ drout = -6.04799226571813 ldrout = 2.64017790273801e-06 wdrout = 5.56320493289501e-06 pdrout = -2.08397656786247e-12
+ pscbe1 = -7045694915.45223 lpscbe1 = 3412.36944588841 wpscbe1 = 5880.58006144451 ppscbe1 = -0.00269507573888488
+ pscbe2 = 1.57248685321277e-07 lpscbe2 = -6.74907666870568e-14 wpscbe2 = -1.13532108438376e-13 ppscbe2 = 5.36712072545703e-20
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.000239280361799599 lalpha0 = -1.06403594001624e-10 walpha0 = -1.18039408524876e-10 palpha0 = 6.32122063994392e-17
+ alpha1 = 0.0
+ beta0 = 167.072591493992 lbeta0 = -5.84147337044429e-05 wbeta0 = -8.43432705373824e-05 pbeta0 = 4.2094322823614e-11
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 6.91148529916801e-07 lagidl = -2.78874550095954e-13 wagidl = -5.3501344157977e-13 pagidl = 2.26010978504906e-19
+ bgidl = -6293856091.45601 lbgidl = 3434.39956040886 wbgidl = 6216.9622148116 pbgidl = -0.00265139494163378
+ cgidl = 12340.278648384 lcgidl = -0.00514934075794066 wcgidl = -0.00923280894801911 pcgidl = 4.12309433654944e-9
+ egidl = 18.5457559325511 legidl = -7.83630041303925e-06 wegidl = -1.3823496115301e-05 pegidl = 6.15539031133483e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -2.12299801008 lkt1 = 6.22465811263969e-07 wkt1 = 1.33324515800914e-06 pkt1 = -5.5480731157535e-13
+ kt2 = -0.019032
+ at = 91051.2130560002 lat = -0.0384669057163777 wat = -0.0492210447867767 pat = 2.33603078558042e-8
+ ute = -3.5531627256832 lute = 1.04979750960925e-06 wute = 1.83102286606809e-06 pute = -8.69003452235916e-13
+ ua1 = 5.52e-10
+ ub1 = -6.91666441205762e-18 lub1 = 2.39533676996255e-24 wub1 = 6.37904740436625e-24 pub1 = -3.02749589811223e-30
+ uc1 = -1.18981061409101e-09 luc1 = 4.04796736038492e-16 wuc1 = 1.12361459408938e-15 puc1 = -4.2090602694588e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 1.81e-6
+ sbref = 1.81e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.72 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 7e-07 wmax = 7.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.893436+0*(0.0/sqrt(l*w*mult))}
+ k1 = 0.57102
+ k2 = 0.0284341
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 180350.0
+ ua = 2.33476787e-9
+ ub = 6.10999999999999e-21
+ uc = -3.2639e-11
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0188609
+ a0 = 0.87668
+ keta = -0.0076977
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.1244
+ b0 = 9.3768e-8
+ b1 = 3.0925e-10
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.10903374+0*(0.009/sqrt(l*w*mult))}
+ nfactor = {1.84191+0*(0.02/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.080000000000001
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.99495
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00129
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 225600350.0
+ pscbe2 = 1.4994384e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.8978653e-5
+ alpha1 = 0.0
+ beta0 = 37.686511
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 3.08e-8
+ bgidl = 1701900000.0
+ cgidl = 1200.0
+ egidl = 1.0890786
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.566
+ kt2 = -0.019032
+ at = 351440.0
+ ute = -1.4104
+ ua1 = 2.2096e-11
+ ub1 = -2.3998e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.73 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 7e-07 wmax = 7.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.881763217933329+0*(0.0/sqrt(l*w*mult))} lvth0 = -2.31991874462181e-7
+ k1 = 0.561944523499999 lk1 = 1.8037146524691e-7
+ k2 = 0.0314860646279499 lk2 = -6.06565761946551e-8
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 246098.9727 lvsat = -1.30673453282342
+ ua = 2.3896607419615e-09 lua = -1.09097387308597e-15
+ ub = -8.37654346666668e-20 lub = 1.78623831382613e-24 wub = 6.88766221184934e-41 pub = 1.40129846432482e-45
+ uc = -2.44562524652332e-11 luc = -1.62628834154475e-16
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0193439410883333 lu0 = -9.60024841418972e-9
+ a0 = 0.856175657168333 la0 = 4.07515612042223e-7
+ keta = -0.00737995988999998 lketa = -6.3149575902062e-9
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.129268878304333 lags = -9.67670087473044e-8
+ b0 = 1.553001244e-07 lb0 = -1.22292635960024e-12
+ b1 = 5.12185004166665e-10 lb1 = -4.03325203381084e-15
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.109922001442166+0*(0.009/sqrt(l*w*mult))} lvoff = 1.76538408584833e-8
+ nfactor = {1.925183895+0*(0.02/sqrt(l*w*mult))} lnfactor = -1.65503535356701e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.32810833333333e-05 lcit = -6.52102188166666e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.080000000000001
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.5930381740625 lpclm = -1.18867632242226e-5
+ pdiblc1 = 0.39
+ pdiblc2 = -0.000119597104030013 lpdiblc2 = 2.80151786037547e-08 ppdiblc2 = 2.52435489670724e-29
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 226179618.700334 lpscbe1 = -11.5127337116428
+ pscbe2 = 1.49915366758833e-08 lpscbe2 = 5.6589427888963e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -1.07243303254001e-05 lalpha0 = 5.90334912398995e-10
+ alpha1 = 0.0
+ beta0 = 36.7986715051499 lbeta0 = 1.7645454824345e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 3.788714e-08 lagidl = -1.40854072644001e-13
+ bgidl = 1821003325.0 lbgidl = -2367.13094304496
+ cgidl = 1068.75666666666 lcgidl = 0.00260840875266669
+ egidl = 0.806343318136665 legidl = 5.61925063292102e-6
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.572562166666668 lkt1 = 1.30420437633331e-7
+ kt2 = -0.019032
+ at = 482913.009166667 lat = -2.61297346798384
+ ute = -1.31478923166666 lute = -1.90022577631766e-06 wute = 3.3881317890172e-21
+ ua1 = 2.2096e-11
+ ub1 = -1.95560693833333e-18 lub1 = -8.82815942340041e-24
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.74 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 7e-07 wmax = 7.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.928454346199995+0*(0.0/sqrt(l*w*mult))} lvth0 = 1.3568208418652e-7
+ k1 = 0.598246429500001 lk1 = -1.05491523740695e-7
+ k2 = 0.0192782061161499 lk2 = 3.54754264423654e-8
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -16896.9181000004 lvsat = 0.764252908870262
+ ua = 2.17008925411549e-09 lua = 6.38063765106081e-16
+ ub = 2.75736303999999e-19 lub = -1.0446940774784e-24
+ uc = -5.71872426042998e-11 luc = 9.51146207946204e-17
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0174117767350001 lu0 = 5.61477300256917e-9
+ a0 = 0.938193028494997 la0 = -2.38338380206728e-7
+ keta = -0.00865092032999998 lketa = 3.69334749061797e-9
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.109793365087 lags = 5.6594867633909e-8
+ b0 = -9.08283732000003e-08 lb0 = 7.15237107600721e-13
+ b1 = -2.99555012500001e-10 lb1 = 2.3588759014325e-15
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1063689556735+0*(0.009/sqrt(l*w*mult))} lvoff = -1.03249733514564e-8
+ nfactor = {1.592088315+0*(0.02/sqrt(l*w*mult))} lnfactor = 9.67959100701005e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.56750000000029e-07 lcit = 3.813865645e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.080000000000001
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.799314522187501 lpclm = 6.95205731766769e-06 wpclm = 4.2351647362715e-22 ppclm = -3.23117426778526e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00551879131209002 lpdiblc2 = -1.63848748178239e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 223862543.898999 lpscbe1 = 6.73330351894037
+ pscbe2 = 1.500292597235e-08 lpscbe2 = -3.30967260673236e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.0001080876029762 lalpha0 = -3.45261537577786e-10
+ alpha1 = 0.0
+ beta0 = 40.3500294845501 lbeta0 = -1.03200687202373e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 9.53857999999984e-09 lagidl = 8.2379497932e-14
+ bgidl = 1344590024.99999 lbgidl = 1384.43322913497
+ cgidl = 1593.73 lcgidl = -0.00152554625799997
+ egidl = 1.93728444559 legidl = -3.28645836932299e-6
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.5463135 lkt1 = -7.62773128999965e-8
+ kt2 = -0.019032
+ at = -42979.0274999999 lat = 1.5282159639515 pat = -1.6940658945086e-21
+ ute = -1.69723230499999 lute = 1.111360448953e-6
+ ua1 = 2.2096e-11
+ ub1 = -3.732379185e-18 lub1 = 5.16321131020101e-24
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.75 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 7e-07 wmax = 7.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.922392946200002+0*(0.0/sqrt(l*w*mult))} lvth0 = 1.12196583746523e-7
+ k1 = 0.581499014000002 lk1 = -4.06019876443979e-8
+ k2 = 0.0220012751288 lk2 = 2.49246232459517e-8
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 313587.194999999 lvsat = -0.516240835747002
+ ua = 2.61870675532099e-09 lua = -1.10014960506475e-15
+ ub = 2.97169768999999e-19 lub = -1.1277401809674e-24 wub = 3.67341984631965e-40 pub = -1.75162308040602e-46
+ uc = -6.06099033194498e-11 luc = 1.08376062001541e-16
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0208186385100001 lu0 = -7.58545363084621e-9
+ a0 = 1.005408782 la0 = -4.98772538737206e-7
+ keta = 0.0199444954899999 lketa = -1.07102450645554e-07 pketa = -5.04870979341448e-29
+ a1 = 0.0
+ a2 = 0.5
+ ags = -0.164308898750999 lags = 1.11863149910062e-6
+ b0 = 3.98057644000001e-08 lb0 = 2.0908207805576e-13
+ b1 = 2.70680104999999e-10 lb1 = 1.49442915167e-16
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.140245475700601+0*(0.009/sqrt(l*w*mult))} lvoff = 1.20932991145546e-7
+ nfactor = {1.68955188500001+0*(0.02/sqrt(l*w*mult))} lnfactor = 5.90326752379012e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.0987460000000008 leta0 = -7.26332516000004e-08 weta0 = -2.11758236813575e-22
+ etab = -0.135611 letab = 2.542163806e-7
+ dsub = 0.788742713016997 ldsub = -8.86286515855669e-07 wdsub = 1.6940658945086e-21
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.830163474460001 lpclm = 6.38481871857286e-7
+ pdiblc1 = 0.243200242714002 lpdiblc1 = 5.6879033958033e-7
+ pdiblc2 = 0.000595784443419997 lpdiblc2 = 2.68980759552488e-9
+ pdiblcb = -0.025
+ drout = 0.685746733930998 ldrout = -4.87218295289055e-07 wdrout = -1.6940658945086e-21
+ pscbe1 = 176358169.740001 lpscbe1 = 190.793751635396
+ pscbe2 = 1.54446788541001e-08 lpscbe2 = -1.74471244169583e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.67672507269e-05 lalpha0 = -6.89237007526466e-11
+ alpha1 = -9.37299999999998e-11 lalpha1 = 3.63166258e-16
+ beta0 = 70.1981777602998 lbeta0 = -0.000125969704029459
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 5.956986112e-08 lagidl = -1.11471703895552e-13
+ bgidl = 2333077820.0 lbgidl = -2445.56158137198
+ cgidl = 759.469000000005 lcgidl = 0.0017068814126
+ egidl = 1.257234475342 legidl = -6.51536754600108e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.489141400000001 lkt1 = -2.9779633156e-7
+ kt2 = -0.019032
+ at = 648226.672 lat = -1.1499296393312
+ ute = -1.37347038 lute = -1.43087505651991e-7
+ ua1 = -4.74957939199999e-10 lua1 = 1.92588519282432e-15 wua1 = -1.97215226305253e-31
+ ub1 = -1.28338197e-18 lub1 = -4.32567329903799e-24
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.76 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 7e-07 wmax = 7.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.886627609400005+0*(0.0/sqrt(l*w*mult))} lvth0 = 4.51508833812392e-8
+ k1 = 0.55984
+ k2 = 0.0361577629399998 lk2 = -1.61312880492397e-9
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 10800.5312000001 lvsat = 0.0513630442124801
+ ua = 2.03203993132e-09 lua = -3.83976792463448e-19
+ ub = -3.25926414000001e-19 lub = 4.03159236844013e-26
+ uc = -2.7970035e-12
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0171172297000001 lu0 = -6.46792675620007e-10
+ a0 = 0.73934
+ keta = -0.0411832982 lketa = 7.48771140572002e-9
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.43242187
+ b0 = 7.5599640000001e-08 lb0 = 1.41982878856e-13
+ b1 = 4.06112019999999e-10 lb1 = -1.04437752692001e-16
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.075734118+0*(0.009/sqrt(l*w*mult))}
+ nfactor = {2.034336336+0*(0.02/sqrt(l*w*mult))} lnfactor = -5.60061794656111e-8
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.0808933194000011 leta0 = -3.916661654724e-8
+ etab = 0.00379637622 letab = -7.11668686201199e-9
+ dsub = 0.31595571
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.1707598
+ pdiblc1 = 0.54661982
+ pdiblc2 = 0.0020306546
+ pdiblcb = -0.025
+ drout = 0.42584153
+ pscbe1 = 278136550.0
+ pscbe2 = 1.4513967e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 3.0
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.056e-10
+ bgidl = 1028500000.0
+ cgidl = 2261.17712399999 lcgidl = -0.0011082206366504
+ egidl = 0.90967406
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.648
+ kt2 = -0.019032
+ at = 38998.0800000001 lat = -0.00786972076799997
+ ute = -1.4498
+ ua1 = 5.524e-10
+ ub1 = -3.5909e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.81e-6
+ sbref = 2.81e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.77 pmos
* DC IV MOS Parameters
+ lmin = 8.0e-07 lmax = 1e-06 wmin = 7e-07 wmax = 7.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.834068679000005+0*(0.0/sqrt(l*w*mult))} lvth0 = -8.17157146602279e-10
+ k1 = 0.55984
+ k2 = 0.0225523675999999 lk2 = 1.02861499594399e-8
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 86976.529000001 lvsat = -0.0152604834634
+ ua = 2.02907384840003e-09 lua = 2.21015932934799e-18
+ ub = 2.24669610000001e-19 lub = -4.41235358905999e-25
+ uc = -2.7970035e-12
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0179542402000001 lu0 = -1.37884205892005e-9
+ a0 = 0.73934
+ keta = -0.032622
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.43242187
+ b0 = 1.04051162e-06 lb0 = -7.01929138852e-13
+ b1 = 1.2537391e-09 lb1 = -8.45772396859999e-16
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.075734118+0*(0.009/sqrt(l*w*mult))}
+ nfactor = {1.91525264000001+0*(0.02/sqrt(l*w*mult))} lnfactor = 4.8144421056003e-8
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.036111000000001
+ etab = -0.0043407
+ dsub = 0.31595571
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.1707598
+ pdiblc1 = 0.54661982
+ pdiblc2 = 0.0020306546
+ pdiblcb = -0.025
+ drout = 0.42584153
+ pscbe1 = 278136550.0
+ pscbe2 = 1.4513967e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 3.0
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -3.47731199999999e-10 lagidl = 3.96483467519999e-16
+ bgidl = 1028500000.0
+ cgidl = 994.06
+ egidl = 0.90967406
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.649686500000001 lkt1 = 1.47501290000162e-9
+ kt2 = -0.019032
+ at = 97460.0000000002 lat = -0.059000516
+ ute = -1.34861000000001 lute = -8.85007740000158e-8
+ ua1 = 5.524e-10
+ ub1 = -3.5909e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.41e-6
+ sbref = 2.41e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.78 pmos
* DC IV MOS Parameters
+ lmin = 6e-07 lmax = 8.0e-07 wmin = 7e-07 wmax = 7.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.014/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.829563443000005+0*(0.0/sqrt(l*w*mult))} lvth0 = -3.85638935220071e-9
+ k1 = 0.534092950000002 lk1 = 1.73689599299996e-8
+ k2 = 0.028832558016 lk2 = 6.04953350480626e-9
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 75470.6066000001 lvsat = -0.00749858821235994
+ ua = 4.584563234107e-09 lua = -1.72172298026859e-15
+ ub = -5.14165594e-18 lub = 3.178887857124e-24 wub = -5.87747175411144e-39 pub = -1.40129846432482e-45
+ uc = -2.68286291190001e-12 luc = -7.69992407322661e-20
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.01806873334 lu0 = -1.45607913116398e-9
+ a0 = 0.570928190000004 la0 = 1.13610607026001e-7
+ keta = 0.0635794199999999 lketa = -6.48974779320003e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = -0.804847112389993 lags = 8.34661655520294e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.000834093863999463+0*(0.009/sqrt(l*w*mult))} lvoff = -5.0527556282146e-8
+ nfactor = {3.73841605999999+0*(0.02/sqrt(l*w*mult))} lnfactor = -1.181761622076e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 2.18649999999999e-05 lcit = -8.00412900000002e-12
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.072247044000001 leta0 = -2.43773752824001e-8
+ etab = -0.0146411811 letab = 6.94870455006e-9
+ dsub = 0.376336362779998 ldsub = -4.07327883653874e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.05547993459999 lpclm = 7.77677971988354e-8
+ pdiblc1 = 0.421065979910004 lpdiblc1 = 8.46986205247131e-8
+ pdiblc2 = -0.0039369499009 lpdiblc2 = 4.02574599630715e-9
+ pdiblcb = -0.025
+ drout = -0.934565625939999 ldrout = 9.17730667397127e-7
+ pscbe1 = -11045416.8499985 lpscbe1 = 195.08215483701
+ pscbe2 = 1.459493376e-08 lpscbe2 = -5.46201762959841e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -8.1316525628e-05 lalpha0 = 5.48561956486488e-11 walpha0 = -5.2194192933043e-26 palpha0 = -3.54194315416888e-32
+ alpha1 = 3.373e-10 lalpha1 = -1.6008258e-16
+ beta0 = -107.343629109 lbeta0 = 7.44378121969314e-05 wbeta0 = -2.71050543121376e-20 pbeta0 = -2.58493941422821e-26
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -6.82447799999999e-08 lagidl = 4.61998325879999e-14 wagidl = 4.41762106923767e-29 pagidl = 3.00926553810506e-36
+ bgidl = -661550600.0 lbgidl = 1140.10813475999
+ cgidl = 1454.56438 lcgidl = -0.000310656254748003
+ egidl = 0.806232427159998 legidl = 6.97817255138621e-8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.751959460000002 lkt1 = 7.04683517159991e-8
+ kt2 = -0.019032
+ at = 10000.0
+ ute = -1.8086978 lute = 2.21874455879997e-7
+ ua1 = 5.53349200000001e-10 lua1 = -6.40330319999736e-19
+ ub1 = -7.6755449e-18 lub1 = 2.75550144954e-24
+ uc1 = -2.80226855999999e-10 luc1 = 1.153747170576e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.02e-6
+ sbref = 2.01e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.79 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 6e-07 wmin = 7e-07 wmax = 7.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.874905510000012+0*(0.0/sqrt(l*w*mult))} lvth0 = 1.76629556460009e-8
+ k1 = 0.714723700000008 lk1 = -6.83583940199973e-8
+ k2 = -0.0634318966079994 lk2 = 4.98382436693568e-8
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 21359.7088000011 lvsat = 0.0181824438835201
+ ua = -2.47267983201399e-09 lua = 1.62764457891244e-15
+ ub = 8.60440408000002e-18 lub = -3.344992228368e-24
+ uc = 5.55978501279998e-12 luc = -3.98895994579486e-18
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0169239913200001 lu0 = -9.12784568472041e-10
+ a0 = 1.28938594 la0 = -2.27369441124001e-7
+ keta = -0.168130592000002 lketa = 4.50720937631996e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.822580059800003 lags = 6.22847195989213e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.137370707712002+0*(0.009/sqrt(l*w*mult))} lvoff = 1.42727206501153e-8
+ nfactor = {-3.15056525999999+0*(0.02/sqrt(l*w*mult))} lnfactor = 2.08774891239599e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -1.37299999999999e-05 lcit = 8.88925800000001e-12
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -0.156355243999999 leta0 = 8.41172706023999e-8
+ etab = 0.0163786358 letab = -7.77330055068001e-9
+ dsub = 0.368580674100002 ldsub = -3.70519385178581e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.89414254160002 lpclm = -3.20261476083356e-7
+ pdiblc1 = 2.16941717718001 lpdiblc1 = -7.45068857699626e-7
+ pdiblc2 = 0.00769304350460004 lpdiblc2 = -1.49384887394316e-9
+ pdiblcb = -0.025
+ drout = 0.995858213260007 ldrout = 1.55151331280068e-9
+ pscbe1 = 400000000.0
+ pscbe2 = 1.35000357480002e-08 lpscbe2 = 4.65018420199242e-16
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 8.98247953940003e-05 lalpha0 = -2.63674753083924e-11
+ alpha1 = 0.0
+ beta0 = 60.2813814380006 lbeta0 = -5.1170178086749e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.37414000000002e-08 lagidl = 7.28919156000005e-15
+ bgidl = 1577749000.00002 lbgidl = 77.3365446000025
+ cgidl = 650.160000000011 lcgidl = 7.11140640000003e-5
+ egidl = 1.04313992120001 legidl = -4.26545711575177e-8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.434910000000002 lkt1 = -8.00033219999992e-8
+ kt2 = -0.019032
+ at = 28730.0 lat = -0.00888925800000001
+ ute = -1.23481360000002 lute = -5.04909854399959e-8
+ ua1 = 5.52e-10
+ ub1 = 1.16016479999997e-18 lub1 = -1.43792637408001e-24
+ uc1 = 2.32853712e-10 luc1 = -1.281333205152e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 1.81e-6
+ sbref = 1.81e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.80 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 4.2e-07 wmax = 7.0e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.822793270985715+0*(0.0/sqrt(l*w*mult))} wvth0 = -5.22612083538525e-8
+ k1 = 0.518816732714286 wk1 = 3.86197683249023e-8
+ k2 = 0.0456003570462571 wk2 = -1.26995282977928e-8
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 432631.854557143 wvsat = -0.186637106873956
+ ua = 3.56563205702014e-09 wua = -9.10588402100754e-16
+ ub = -1.41482221072857e-18 wub = 1.05119996576815e-24
+ uc = -1.77404223410429e-11 wuc = -1.10219081577859e-17
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0195344485918857 wu0 = -4.98288554082683e-10
+ a0 = 0.831242302428572 wa0 = 3.36146269125523e-8
+ keta = -0.0134352972285714 wketa = 4.24465147930823e-9
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.151636820703 wags = -2.01496910087966e-8
+ b0 = 2.08948540128571e-07 wb0 = -8.52101028649566e-14
+ b1 = -8.99767160714285e-10 wb1 = 8.94426059427785e-16
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0874468104385716+0*(0.009/sqrt(l*w*mult))} wvoff = -1.59699241418266e-8
+ nfactor = {1.89940092128572+0*(0.02/sqrt(l*w*mult))} wnfactor = -4.2531553603486e-8
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 2.62704125588647e-05 wcit = -1.20367861293979e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.080000000000001
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.49161676991071 wpclm = -1.10722808971287e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00129
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 226586201.887857 wpscbe1 = -0.729329283229163
+ pscbe2 = 1.49851618059429e-08 wpscbe2 = 6.82254227469533e-18
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 5.01438771256714e-05 walpha0 = -2.30559081472752e-11
+ alpha1 = -1.64212857142857e-10 walpha1 = 1.21484014862857e-16
+ beta0 = 94.6462217562714 wbeta0 = -4.21385661786466e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 6.49562742857143e-08 wagidl = -2.52686750914743e-14
+ bgidl = 2450053777.14286 wbgidl = -553.481171715177
+ cgidl = 871.574285714287 wcgidl = 0.000242968029725714
+ egidl = -0.406771457265713 wegidl = 1.10662388896495e-6
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.582864660428572 wkt1 = 1.24764083264153e-8
+ kt2 = -0.019032
+ at = 851698.048 wat = -0.370088902878208
+ ute = -1.35391077714286 wute = -4.1790501112823e-8
+ ua1 = -1.10188189051428e-09 wua1 = 8.31514347490906e-16
+ ub1 = -1.17608578857143e-18 wub1 = -9.0529887875801e-25
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.81 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 4.2e-07 wmax = 7.0e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.784469480177342+0*(0.0/sqrt(l*w*mult))} lvth0 = -7.61670012800078e-07 wvth0 = -7.19775180169314e-08 pvth0 = 3.91853768029828e-13
+ k1 = 0.44367408227146 lk1 = 1.49343012049099e-06 wk1 = 8.74959993391094e-08 pk1 = -9.71395540914958e-13
+ k2 = 0.0693006152681457 lk2 = -4.71033152056747e-07 wk2 = -2.79750533054143e-08 pk2 = 3.03594949316473e-13
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 663932.384915116 lvsat = -4.59700552065257 wvsat = -0.309111487023094 pvsat = 2.43412931571205e-6
+ ua = 4.38821426168721e-09 lua = -1.63484922848761e-14 wua = -1.478521899679e-15 pua = 1.12874510909687e-20
+ ub = -2.36279072994451e-18 lub = 1.88404951320092e-23 wub = 1.68601379734537e-24 pub = -1.26166709770645e-29
+ uc = 1.48339518889436e-11 luc = -6.47402658071288e-16 wuc = -2.90667360204026e-17 puc = 3.58633735838364e-22
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0226290212940561 lu0 = -6.15033946265561e-08 wu0 = -2.43028919587291e-09 pu0 = 3.83977399553239e-14
+ a0 = 0.750827823849432 la0 = 1.59820559596895e-06 wa0 = 7.79359056979899e-08 pa0 = -8.80867687349049e-13
+ keta = -0.0136185297032398 lketa = 3.64167214104462e-09 wketa = 4.61526899355557e-09 pketa = -7.36587484866029e-15
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.176673816467263 lags = -4.97600276016418e-07 wags = -3.50699836331826e-08 pags = 2.96534847792622e-13
+ b0 = 4.14870467792657e-07 lb0 = -4.09261594355264e-12 wb0 = -1.92029101760514e-13 pb0 = 2.12298487544965e-18
+ b1 = 7.8672947324212e-08 lb1 = -1.58147587130212e-12 wb1 = -5.78230193213203e-14 pb1 = 1.16698573996422e-18
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0951575232209244+0*(0.009/sqrt(l*w*mult))} lvoff = 1.53247332264152e-07 wvoff = -1.09227019301622e-08 pvoff = -1.00311522567947e-13
+ nfactor = {2.08322493862473+0*(0.02/sqrt(l*w*mult))} lnfactor = -3.65342881500602e-06 wnfactor = -1.16918131909401e-07 pnfactor = 1.47840348919874e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 3.75344314434153e-05 lcit = -2.2386786972289e-10 wcit = -1.79425299184462e-11 pcit = 1.1737429550982e-16
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.080000000000001
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 4.07184235343675 lpclm = -3.14063513823466e-05 wpclm = -1.83380941668436e-06 ppclm = 1.44405132410276e-11
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00225565206719492 lpdiblc2 = -1.91919485746721e-08 wpdiblc2 = -1.75719983587551e-09 ppdiblc2 = 3.49236438580914e-14
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 228116704.271542 lpscbe1 = -30.418122674786 wpscbe1 = -1.43304815723798 ppscbe1 = 1.39861311333755e-5
+ pscbe2 = 1.49776388095421e-08 lpscbe2 = 1.49516544266633e-16 wpscbe2 = 1.02815859277797e-17 ppscbe2 = -6.8747108987616e-23
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -2.83352237750343e-05 lalpha0 = 1.55974073876117e-09 walpha0 = 1.30284685304657e-11 palpha0 = -7.17162552719429e-16
+ alpha1 = -1.64212857142857e-10 walpha1 = 1.21484014862857e-16
+ beta0 = 92.3004356600855 lbeta0 = 4.6621560347256e-05 wbeta0 = -4.10599831147647e-05 pbeta0 = -2.1436406961427e-11
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.48336937612286e-07 lagidl = -1.65715733135028e-12 wagidl = -8.17103184743785e-14 pagidl = 1.12175508557787e-18
+ bgidl = 2822606772.85486 lbgidl = -7404.34176857771 wbgidl = -740.982224309232 pbgidl = 0.0037265084198858
+ cgidl = 616.407856582143 lcgidl = 0.00507133071242969 wcgidl = 0.00033464584030529 pcgidl = -1.82205981414485e-9
+ egidl = -1.15379442362774 legidl = 1.48467826472587e-05 wegidl = 1.45010206080634e-06 pegidl = -6.82649127407895e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.589717776972331 lkt1 = 1.36202950060603e-07 wkt1 = 1.26916518816893e-08 pkt1 = -4.27787956364434e-15
+ kt2 = -0.019032
+ at = 1311448.7258984 lat = -9.13736082295953 wat = -0.612947409095269 pat = 4.8267156676616e-6
+ ute = -1.22123083928362 lute = -2.63696069297722e-06 wute = -6.9214124451409e-08 pute = 5.45033544405065e-13
+ ua1 = -1.8394549152346e-09 lua1 = 1.46589688371064e-14 wua1 = 1.3771679208869e-15 pua1 = -1.0844646509816e-20
+ ub1 = 7.11289338715214e-20 lub1 = -2.47878937226647e-23 wub1 = -1.49937109131366e-24 pub1 = 1.18069475956586e-29
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.82 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 4.2e-07 wmax = 7.0e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.927404754024259+0*(0.0/sqrt(l*w*mult))} lvth0 = 3.6388809463486e-07 wvth0 = -7.76484093243811e-10 pvth0 = -1.6882589370564e-13
+ k1 = 0.72461608968835 lk1 = -7.18875811114052e-07 wk1 = -9.34877691287005e-08 pk1 = 4.53779242261657e-13
+ k2 = -0.024242421961623 lk2 = 2.6558084891279e-07 wk2 = 3.21963865694242e-08 pk2 = -1.7023107112193e-13
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -112526.666283743 lvsat = 1.51729892391796 wvsat = 0.0707465051873402 pvsat = -5.57100429748229e-7
+ ua = 1.94071927846393e-09 lua = 2.92455171001393e-15 wua = 1.69686990507129e-16 pua = -1.69153463569105e-21
+ ub = 7.94382329725916e-19 lub = -6.02097984367158e-24 wub = -3.8369225524793e-25 pub = 3.68143630468665e-30
+ uc = -9.27885673824173e-11 luc = 2.0008163218297e-16 wuc = 2.63377176655521e-17 puc = -7.76541751570553e-23
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0139735272299217 lu0 = 6.65515893087676e-09 wu0 = 2.5436032308589e-09 pu0 = -7.69673348218332e-16
+ a0 = 0.922408114394596 la0 = 2.47079440042011e-07 wa0 = 1.16776163118224e-08 pa0 = -3.59110161748735e-13
+ keta = -0.0142473534210017 lketa = 8.59340738893238e-09 wketa = 4.14021881499071e-09 pketa = -3.62504471253339e-15
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.0877004526207974 lags = 2.03029374928958e-07 wags = 1.63442482708468e-08 pags = -1.08331662758848e-13
+ b0 = -3.40478239683078e-07 lb0 = 1.85545298833579e-12 wb0 = 1.84689972624716e-13 pb0 = -8.4352714770428e-19
+ b1 = -2.30344592768913e-07 lb1 = 8.51913649915206e-13 wb1 = 1.70186398752043e-13 pb1 = -6.28497223596294e-19
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.109462157006333+0*(0.009/sqrt(l*w*mult))} lvoff = 2.65890601470734e-07 wvoff = 2.28833797322477e-09 pvoff = -2.04343177391157e-13
+ nfactor = {0.454955077970071+0*(0.02/sqrt(l*w*mult))} lnfactor = 9.16854502970516e-06 wnfactor = 8.41246620221792e-07 pnfactor = -6.06676066793356e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 2.85451826785714e-07 lcit = 6.94529451662218e-11 wcit = -9.52130966487643e-14 pcit = -2.3166185535106e-17
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.080000000000001
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.320256395028067 lpclm = 3.17966942231443e-06 wpclm = -3.5440528624004e-07 ppclm = 2.79079747543076e-12
+ pdiblc1 = 0.39
+ pdiblc2 = -0.00160695620158476 lpdiblc2 = 1.12245464986603e-08 wpdiblc2 = 5.27159950762653e-09 ppdiblc2 = -2.04253394522497e-14
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 221996985.269693 lpscbe1 = 17.7722165771775 wpscbe1 = 1.38013281172687 ppscbe1 = -8.16654372483511e-6
+ pscbe2 = 1.50077482922714e-08 lpscbe2 = -8.75835884335028e-17 wpscbe2 = -3.56753298857097e-18 ppscbe2 = 4.03091628310828e-23
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.000320671300668863 lalpha0 = -1.18854603862475e-09 walpha0 = -1.57268569218241e-10 palpha0 = 6.23858500736538e-16
+ alpha1 = -3.23277641214286e-10 lalpha1 = 1.25257154864887e-15 walpha1 = 2.39159505859764e-16 palpha1 = -9.2664742140424e-22
+ beta0 = 155.707729316783 lbeta0 = -0.00045268551428177 wbeta0 = -8.53411649050863e-05 pbeta0 = 3.2726018716464e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -9.97679266476428e-08 lagidl = 2.96569232750957e-13 wagidl = 8.08645163918996e-14 pagidl = -1.58456709060125e-19
+ bgidl = 1872799260.50415 lbgidl = 75.0124681791567 wbgidl = -390.767079589029 pbgidl = 0.000968704241272093
+ cgidl = 1318.94400496786 lcgidl = -0.000460860441648461 wcgidl = 0.000203285579980799 pcgidl = -7.87650308193604e-10
+ egidl = 0.767235038530006 legidl = -2.80555955448688e-07 wegidl = 8.65597871145357e-07 pegidl = -2.22375458217457e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.578641264121429 lkt1 = 4.89798419648882e-08 wkt1 = 2.39159505859765e-08 pkt1 = -9.26647421404239e-14
+ kt2 = -0.019032
+ at = -252610.506427736 lat = 3.17898000791585 wat = 0.155084529584823 pat = -1.22122863666865e-6
+ ute = -1.74813303590286 lute = 1.51218334452063e-06 wute = 3.765615711901e-08 pute = -2.96527174849356e-13
+ ua1 = 2.2096e-11
+ ub1 = -3.732379185e-18 lub1 = 5.163211310201e-24
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.83 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 4.2e-07 wmax = 7.0e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.898762048531878+0*(0.0/sqrt(l*w*mult))} lvth0 = 2.52909067934079e-07 wvth0 = -1.74820435712861e-08 pvth0 = -1.0409853295202e-13
+ k1 = 0.568183535316714 lk1 = -1.12762235945712e-07 wk1 = 9.85073786798031e-09 pk1 = 5.33838630523173e-14
+ k2 = 0.0261282076142353 lk2 = 7.04148075581689e-08 wk2 = -3.05308814499511e-09 pk2 = -3.36534563934412e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 647450.524108985 lvsat = -1.4273086979777 wvsat = -0.246990755421511 pvsat = 6.74004360206826e-7
+ ua = 3.2054282874797e-09 lua = -1.97568981631857e-15 wua = -4.34054242604876e-16 pua = 6.4772114612473e-22
+ ub = 4.9475512345712e-19 lub = -4.86004427026252e-24 wub = -1.46172854885961e-25 pub = 2.76114363604417e-30
+ uc = -9.04878065320654e-11 luc = 1.91167104192197e-16 wuc = 2.210355328508e-17 puc = -6.12484818484783e-23
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0214149990651467 lu0 = -2.2177567841886e-08 wu0 = -4.41185153255299e-10 pu0 = 1.07951877248705e-14
+ a0 = 1.43403682373026 la0 = -1.73527715714994e-06 wa0 = -3.17097310759877e-07 pa0 = 9.14761170683272e-13
+ keta = 0.0549401372757495 lketa = -2.594804440647e-07 wketa = -2.58896358105304e-08 pketa = 1.12728630019511e-13
+ a1 = 0.0
+ a2 = 0.5
+ ags = -0.645545053372945 lags = 3.04406241245231e-06 wags = 3.56016582244697e-07 pags = -1.42442608797393e-12
+ b0 = -2.71364622102429e-09 lb0 = 5.46750294507712e-13 wb0 = 3.14556898997913e-14 pb0 = -2.49805595858288e-19
+ b1 = 7.75892964202037e-08 lb1 = -3.41206997136946e-13 wb1 = -5.72000030755225e-14 pb1 = 2.52534128924793e-19
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.120178083575282+0*(0.009/sqrt(l*w*mult))} lvoff = 3.07410530554781e-07 wvoff = -1.4845776424742e-08 pvoff = -1.37955337744795e-13
+ nfactor = {2.5001784747307+0*(0.02/sqrt(l*w*mult))} lnfactor = 1.24412245661642e-06 wnfactor = -5.99698308576412e-07 pnfactor = -4.83675446812033e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.82106428571429e-05 wcit = -6.07420074314286e-12
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.7605878573 leta0 = -2.63700571189458e-06 weta0 = -4.89627958663111e-07 peta0 = 1.89711248863609e-12
+ etab = -1.761741051715 letab = 6.55481987897494e-06 wetab = 1.20300450773855e-06 petab = -4.66116126568379e-12
+ dsub = 0.702617524568302 ldsub = -5.52585860692343e-07 wdsub = 6.37150699135931e-08 pdsub = -2.46870409887208e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.952603559599785 lpclm = -1.75215375788665e-06 wpclm = -9.05806852260728e-08 ppclm = 1.76858267634204e-12
+ pdiblc1 = 0.299820890564371 lpdiblc1 = 3.4940797741929e-07 wpdiblc1 = -4.18877287971127e-08 ppdiblc1 = 1.62298193997292e-13
+ pdiblc2 = -0.000544206756770204 lpdiblc2 = 7.10681749978184e-09 wpdiblc2 = 8.43360929935914e-10 ppdiblc2 = -3.26768625912969e-15
+ pdiblcb = -0.025
+ drout = 0.507881521591337 ldrout = 2.01938256442206e-07 wdrout = 1.31583972628033e-07 pdrout = -5.09835260344578e-13
+ pscbe1 = 200894961.755213 lpscbe1 = 99.5341168863779 wpscbe1 = -18.152220585687 ppscbe1 = 6.75135127487844e-5
+ pscbe2 = 1.57772737592556e-08 lpscbe2 = -3.06918696281048e-15 wpscbe2 = -2.46052380454478e-16 ppscbe2 = 9.79840952822492e-22
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.58432893087974e-05 lalpha0 = -8.49514258090363e-11 walpha0 = 6.83542961266642e-13 palpha0 = 1.18572468858168e-17
+ alpha1 = -2.47646711e-10 lalpha1 = 9.595319464406e-16 walpha1 = 1.13866967130956e-16 palpha1 = -4.41188950845602e-22
+ beta0 = 122.167933077863 lbeta0 = -0.000322732219774453 wbeta0 = -3.84470171049119e-05 pbeta0 = 1.45564122098084e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 6.0329560900184e-08 lagidl = -3.23744492501853e-13 wagidl = -5.62022858581014e-16 pagidl = 1.57038559919787e-19
+ bgidl = 3533512364.81443 lbgidl = -6359.58652578147 wbgidl = -888.076674515538 pbgidl = 0.00289557999777435
+ cgidl = -37.8195629799984 lcgidl = 0.00479605567872231 wcgidl = 0.000589830889738352 pcgidl = -2.28535876538022e-9
+ egidl = 1.36526190716076 legidl = -2.59767086064543e-06 wegidl = -7.99182619497958e-08 pegidl = 1.4397422271159e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.3967913734 lkt1 = -6.55615744624359e-07 wkt1 = -6.83201802785734e-08 pkt1 = 2.64713370507361e-13
+ kt2 = -0.019032
+ at = 1297133.36266747 lat = -2.82565758728044 wat = -0.480058574129033 pat = 1.23969683298106e-6
+ ute = -1.11806004061629 lute = -9.29097483016707e-07 wute = -1.88951547434713e-07 pute = 5.81487037214502e-13
+ ua1 = -4.749579392e-10 lua1 = 1.92588519282432e-15 wua1 = 6.16297582203915e-33 pua1 = 1.17549435082229e-38
+ ub1 = -6.87262548297003e-19 lub1 = -6.63539761036844e-24 wub1 = -4.41006763698192e-25 pub1 = 1.70872480662502e-30
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.84 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 4.2e-07 wmax = 7.0e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.014/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.759630979567135+0*(0.0/sqrt(l*w*mult))} lvth0 = -7.90603394722988e-09 wvth0 = -9.39515987638342e-08 pvth0 = 3.92512952119325e-14
+ k1 = 0.495082918253468 lk1 = 2.42721808010503e-08 wk1 = 4.79070300477579e-08 pk1 = -1.79564622678939e-14
+ k2 = 0.0763329512751107 lk2 = -2.36990049085081e-08 wk2 = -2.97214436295616e-08 pk2 = 1.63390427979271e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -245628.445496926 lvsat = 0.246857138445537 wvsat = 0.189705131244479 pvsat = -1.44625748937239e-7
+ ua = 1.87080534224814e-09 lua = 5.26194356812522e-16 wua = 1.19280704057009e-16 pua = -3.8956054488764e-22
+ ub = -2.14879000544918e-18 lub = 9.55454283852367e-26 wub = 1.34854719349974e-24 pub = -4.08585666596602e-32
+ uc = 2.18321427016865e-11 luc = -1.93878726413948e-17 wuc = -1.82205438434229e-17 puc = 1.43430706286133e-23
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.00811605659368213 lu0 = 2.75262971512148e-09 wu0 = 6.65903185936153e-09 pu0 = -2.514879086981e-15
+ a0 = 0.154157581940106 la0 = 6.63984469509876e-07 wa0 = 4.32915612151037e-07 pa0 = -4.91213054605529e-13
+ keta = -0.0991959401084917 lketa = 2.94630465997985e-08 wketa = 4.29175204333345e-08 pketa = -1.62572650752385e-14
+ a1 = 0.0
+ a2 = 0.5
+ ags = 1.01869460436079 lags = -7.57212499353375e-08 wags = -4.33722223789172e-07 pags = 5.60182778171629e-14
+ b0 = 7.99356689979572e-08 lb0 = 3.91815888198209e-13 wb0 = -3.20777690857277e-15 pb0 = -1.84825460979329e-19
+ b1 = -1.9466398691831e-07 lb1 = 1.69159007809431e-13 wb1 = 1.44312078914166e-13 pb1 = -1.25220419973077e-19
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {0.083199625119854+0*(0.009/sqrt(l*w*mult))} lvoff = -7.38413221651207e-08 wvoff = -1.17578547425096e-07 pvoff = 5.46275147724676e-14
+ nfactor = {3.82930681900451+0*(0.02/sqrt(l*w*mult))} lnfactor = -1.24746153755926e-06 wnfactor = -1.32791198344481e-06 pnfactor = 8.81433908096259e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.82106428571429e-05 wcit = -6.07420074314286e-12
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -0.88183026575019 leta0 = 4.41871301575309e-07 weta0 = 7.12219057399771e-07 peta0 = -3.55869927675389e-13
+ etab = 3.26118111992112 letab = -2.86115002397413e-06 wetab = -2.40980020385111e-06 petab = 2.1114024466622e-12
+ dsub = 0.419783713059409 ldsub = -2.23855976377726e-08 wdsub = -7.68115413513387e-08 pdsub = 1.65607755900337e-14
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -1.27463339863186 lpclm = 2.4230246440144e-06 wpclm = 1.80909210677506e-06 ppclm = -1.79254393954328e-12
+ pdiblc1 = 0.252364866089742 lpdiblc1 = 4.38369040899431e-07 wpdiblc1 = 2.17688637882994e-07 ppdiblc1 = -3.24303662981235e-13
+ pdiblc2 = 0.00307826986520225 lpdiblc2 = 3.16122824232268e-10 wpdiblc2 = -7.75021582735567e-10 ppdiblc2 = -2.33866400875734e-16
+ pdiblcb = -0.025
+ drout = 1.42797821529972 ldrout = -1.52287500558353e-06 wdrout = -7.41376711237993e-07 pdrout = 1.12661683763068e-12
+ pscbe1 = 277170835.433002 lpscbe1 = -43.4526359100046 wpscbe1 = 0.714431773806609 ppscbe1 = 3.21460862356777e-5
+ pscbe2 = 1.43440492679962e-08 lpscbe2 = -3.82464331495614e-16 wpscbe2 = 1.25704458465491e-16 ppscbe2 = 2.82945582583135e-22
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -2.63080772516525e-06 lalpha0 = -1.282788350917e-11 walpha0 = 1.94633501144635e-12 palpha0 = 9.49001690854994e-18
+ alpha1 = 2.64212857142857e-10 walpha1 = -1.21484014862857e-16
+ beta0 = -42.8979873509509 lbeta0 = -1.32996453385983e-05 wbeta0 = 3.39551474502841e-05 pbeta0 = 9.83902442291363e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -1.39084436286286e-07 lagidl = 5.00769866239032e-14 wagidl = 1.02972232084449e-13 pagidl = -3.70467543964171e-20
+ bgidl = 451117977.291107 lbgidl = -581.330006930237 wbgidl = 427.144910871949 pbgidl = 0.000430065613806962
+ cgidl = 3864.28531151251 lcgidl = -0.00251883011900136 wcgidl = -0.00118597302468901 pcgidl = 1.04356325260531e-9
+ egidl = -1.04356725754166 legidl = 1.91792029150574e-06 wegidl = 1.44500011375205e-06 pegidl = -1.41886975997478e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.821210408011429 lkt1 = 1.40000177658224e-07 wkt1 = 1.28140367005223e-07 pkt1 = -1.03571571430844e-13
+ kt2 = -0.019032
+ at = -449013.498595428 lat = 0.44766931884299 wat = 0.361029013798583 pat = -3.37005959348052e-7
+ ute = -1.757017755156 lute = 2.68692648659437e-07 wute = 2.27278466393388e-07 pute = -1.98777746707657e-13
+ ua1 = 5.524e-10
+ ub1 = -3.78497591764886e-18 lub1 = -8.28424128181451e-25 wub1 = 1.43576587572953e-25 pub1 = 6.12864856332126e-31
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.81e-6
+ sbref = 2.81e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.85 pmos
* DC IV MOS Parameters
+ lmin = 8.0e-07 lmax = 1e-06 wmin = 4.2e-07 wmax = 7.0e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.02/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.547696988363743+0*(0.0/sqrt(l*w*mult))} lvth0 = -1.93263502653715e-07 wvth0 = -2.11856631245941e-07 pvth0 = 1.42371036620783e-13
+ k1 = 0.20871570995822 lk1 = 2.74728941176073e-07 wk1 = 2.59760345275748e-07 pk1 = -2.03243371766293e-13
+ k2 = 0.14962794730278 lk2 = -8.78028084343076e-08 wk2 = -9.40100055617977e-08 pk2 = 7.25658190638609e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -35442.6009042426 lvsat = 0.0630285987647762 wvsat = 0.090565182626639 pvsat = -5.79179498760759e-8
+ ua = 1.37869059723412e-09 lua = 9.56597912801786e-16 wua = 4.81150927679518e-16 pua = -7.06052242467885e-22
+ ub = -2.08492703438293e-18 lub = 3.96908738906989e-26 wub = 1.70863035912792e-24 pub = -3.55787303318067e-31
+ uc = -6.64839115328354e-13 luc = 2.87987655766459e-19 wuc = -1.57736668312255e-18 puc = -2.13052115785404e-25
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.00439496485741656 lu0 = 6.00709654765938e-09 wu0 = 1.00310976613418e-08 pu0 = -5.46408783739298e-15
+ a0 = 1.64395242732151 la0 = -6.38990102260697e-07 wa0 = -6.69228655282742e-07 pa0 = 4.72722321692055e-13
+ keta = -0.159840661881006 lketa = 8.25029202620394e-08 wketa = 9.41158571849206e-08 pketa = -6.10353303981757e-14
+ a1 = 0.0
+ a2 = 0.5
+ ags = 2.47098540524049 lags = -1.34589478438473e-06 wags = -1.50812114911677e-06 pags = 9.95687577908685e-13
+ b0 = 2.30863812151911e-06 lb0 = -1.55740727677679e-12 wb0 = -9.38154913317832e-13 pb0 = 6.3287930452421e-19
+ b1 = -5.47057574661141e-09 lb1 = 3.69045039866406e-15 wb1 = 4.97462122626374e-15 pb1 = -3.35587947923752e-21
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {0.0598655528661675+0*(0.009/sqrt(l*w*mult))} lvoff = -5.34333425720465e-08 wvoff = -1.00316094108107e-07 pvoff = 3.95297731014297e-14
+ nfactor = {5.06015459047505+0*(0.02/sqrt(l*w*mult))} lnfactor = -2.3239609984874e-06 wnfactor = -2.32658588335364e-06 pnfactor = 1.75487410095653e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.82106428571428e-05 wcit = -6.07420074314286e-12
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.745355985715997 leta0 = -9.81265793957019e-07 weta0 = -5.24696603452751e-07 peta0 = 7.25936509306227e-13
+ etab = -0.00595581767477444 letab = -3.71205835276187e-09 wetab = 1.19485759532743e-09 petab = 2.74616592113983e-15
+ dsub = 1.50686075041892 ldsub = -9.73143174512402e-07 wdsub = -8.81026785281757e-07 pdsub = 7.19927427931578e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.61741297744064 lpclm = -1.06359116498617e-07 wpclm = -3.30432234057881e-07 ppclm = 7.86840489492102e-14
+ pdiblc1 = 0.648793585835858 lpdiblc1 = 9.16524826094755e-08 wpdiblc1 = -7.5587743270305e-08 ppdiblc1 = -6.78041400245594e-14
+ pdiblc2 = 0.0329018424124245 lpdiblc2 = -2.57675737255683e-08 wpdiblc2 = -2.28383812588804e-08 ppdiblc2 = 1.90627479718806e-14
+ pdiblcb = -0.025
+ drout = -2.33548106260975 ldrout = 1.76864647887609e-06 wdrout = 2.04281540872232e-06 pdrout = -1.30843759048662e-12
+ pscbe1 = 227113593.710494 lpscbe1 = 0.32742770050163 wpscbe1 = 37.7465789711514 ppscbe1 = -2.4222970311993e-7
+ pscbe2 = 1.14529870164302e-08 lpscbe2 = 2.14605871372399e-15 wpscbe2 = 2.26450074792499e-15 ppscbe2 = -1.58764565217815e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -7.56442770279975e-05 lalpha0 = 5.10296967430871e-11 walpha0 = 5.59614075478045e-11 palpha0 = -3.77515655317489e-17
+ alpha1 = 8.18102824285712e-10 lalpha1 = -4.84432165263141e-16 walpha1 = -5.31249596995273e-16 palpha1 = 3.58380978133011e-22
+ beta0 = -264.210125378699 lbeta0 = 0.00018025995058047 wbeta0 = 0.00019768098191466 pbeta0 = -1.3335559039963e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 3.41977497310129e-06 lagidl = -3.06250145282647e-12 wagidl = -2.53019309615128e-12 pagidl = 2.26591964167855e-18
+ bgidl = -1266898347.62541 lbgidl = 921.247070841741 wbgidl = 1698.12651597988 pbgidl = -0.000681534898020438
+ cgidl = 27284.1091761628 lcgidl = -0.0230018080710245 wcgidl = -0.0194492732203285 pcgidl = 1.70166456037116e-8
+ egidl = 7.99695722673503 legidl = -5.98892242244266e-06 wegidl = -5.24314373761791e-06 pegidl = 4.43058085243339e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.5409677358 lkt1 = -1.05100063457891e-07 wkt1 = -8.04297068801029e-08 pkt1 = 7.88438151892618e-14
+ kt2 = -0.019032
+ at = 241080.564857142 lat = -0.155886949052628 wat = -0.106249919399055 pat = 7.16761956266022e-8
+ ute = -1.34861 lute = -8.85007740000006e-8
+ ua1 = 5.524e-10
+ ub1 = -4.73217935714285e-18 wub1 = 8.44313903296857e-25
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.41e-6
+ sbref = 2.41e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.86 pmos
* DC IV MOS Parameters
+ lmin = 6e-07 lmax = 8.0e-07 wmin = 4.2e-07 wmax = 7.0e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.02/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.847818606783395+0*(0.0/sqrt(l*w*mult))} lvth0 = 9.19854113218156e-09 wvth0 = 1.35050971463001e-08 pvth0 = -9.65798535262321e-15
+ k1 = 0.582278497340552 lk1 = 2.27234848079524e-08 wk1 = -3.56474751803516e-08 pk1 = -3.96125608660945e-15
+ k2 = 0.0114629563233974 lk2 = 5.4032944803838e-09 wk2 = 1.28499618537806e-08 pk2 = 4.78085045311753e-16
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 107237.844939003 lvsat = -0.0332236300010769 wvsat = -0.0235012758542408 pvsat = 1.90312830151256e-8
+ ua = 8.00610106472075e-09 lua = -3.5142531885647e-15 wua = -2.53124000093673e-15 pua = 1.32610667797663e-21
+ ub = -1.21545663850246e-17 lub = 6.83266957983359e-24 wub = 5.18812309558745e-24 pub = -2.70305310333367e-30
+ uc = -1.12648625243293e-12 luc = 5.99414814457212e-19 wuc = -1.1514012271671e-18 puc = -5.00408412372952e-25
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0149538312600317 lu0 = -1.11591472754484e-09 wu0 = 2.30439209915219e-09 pu0 = -2.51652265139834e-16
+ a0 = -0.261997185557855 la0 = 6.4676350658772e-07 wa0 = 6.161948611362e-07 pa0 = -3.94424382484163e-13
+ keta = 0.257880452987162 lketa = -1.99291743828026e-07 wketa = -1.4374312699977e-07 pketa = 9.94243403328167e-14
+ a1 = 0.0
+ a2 = 0.5
+ ags = -2.69000097647244 lags = 2.13570662871881e-06 wags = 1.39462928803273e-06 pags = -9.62507866992373e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {0.173541613355992+0*(0.009/sqrt(l*w*mult))} lvoff = -1.30119212978482e-07 wvoff = -1.29002450698521e-07 pvoff = 5.88815892573228e-14
+ nfactor = {2.96722258021198+0*(0.02/sqrt(l*w*mult))} lnfactor = -9.12069064363933e-07 wnfactor = 5.70525851573251e-07 pnfactor = -1.99517475425156e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 6.90433538571429e-05 lcit = -3.42917468406e-11 wcit = -3.49023574700988e-11 pcit = 1.94474745280045e-17
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -2.15510580541483 leta0 = 9.75385730339837e-07 weta0 = 1.64778672858569e-06 peta0 = -7.39620746486908e-13
+ etab = -0.178528044650714 letab = 1.12705165965207e-07 wetab = 1.21242846107364e-07 petab = -7.82382071290799e-14
+ dsub = -0.458061590457637 ldsub = 3.52393436642924e-07 wdsub = 6.17284268213391e-07 pdsub = -2.90833208756249e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.56423572956765 lpclm = -7.0485745083491e-08 wpclm = -3.76375502093887e-07 ppclm = 1.096773775663e-13
+ pdiblc1 = 0.267681264803853 lpdiblc1 = 3.48750854377667e-07 wpdiblc1 = 1.13473398696667e-07 ppdiblc1 = -1.95344786395479e-13
+ pdiblc2 = -0.0337336072400407 lpdiblc2 = 1.91847006099847e-08 wpdiblc2 = 2.2043447912867e-08 ppdiblc2 = -1.12145339873802e-14
+ pdiblcb = -0.025
+ drout = -2.50090581321865 ldrout = 1.88024201563686e-06 wdrout = 1.158772205188e-06 pdrout = -7.1206204538236e-13
+ pscbe1 = -239924854.762699 lpscbe1 = 315.391565040517 wpscbe1 = 169.324092650063 ppscbe1 = -8.90044204309134e-5
+ pscbe2 = 1.23698784356822e-08 lpscbe2 = 1.52752376229657e-15 wpscbe2 = 1.64608702870897e-15 ppscbe2 = -1.17046375719503e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -0.000137503834312634 lalpha0 = 9.27601540873029e-11 walpha0 = 4.15671462156575e-11 palpha0 = -2.80411968370825e-17
+ alpha1 = 3.373e-10 lalpha1 = -1.6008258e-16
+ beta0 = -124.530100342513 lbeta0 = 8.60318056910592e-05 wbeta0 = 1.27144826726679e-05 pbeta0 = -8.57719001098178e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -3.64831493087171e-06 lagidl = 1.70563199639371e-12 wagidl = 2.64852157733429e-12 pagidl = -1.22764127705481e-18
+ bgidl = -4419883130.64946 lbgidl = 3048.25060546977 wbgidl = 2780.39937284435 pbgidl = -0.00141163616726121
+ cgidl = -20559.7383709054 lcgidl = 0.00927365148422771 wcgidl = 0.0162860931179088 pcgidl = -7.09043252806328e-9
+ egidl = -3.72969645874728 legidl = 1.92187815378371e-06 wegidl = 3.35566204607866e-06 pegidl = -1.37017352924832e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.918126450142857 lkt1 = 1.493312052378e-07 wkt1 = 1.22929674639725e-07 pkt1 = -5.83424235840133e-14
+ kt2 = -0.019032
+ at = 10000.0
+ ute = -1.41902069 lute = -4.10017225259992e-08 wute = -2.8828156726956e-07 pute = 1.94474745280045e-13
+ ua1 = 5.533492e-10 lua1 = -6.40330320000131e-19
+ ub1 = -1.15250801716429e-17 lub1 = 4.5824908894617e-24 wub1 = 2.8478707958203e-24 pub1 = -1.35159947969631e-30
+ uc1 = -5.610749427192e-10 luc1 = 3.04834836358372e-16 wuc1 = 2.07770291162517e-16 puc1 = -1.40161838418234e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.02e-6
+ sbref = 2.01e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.87 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 6e-07 wmin = 4.2e-07 wmax = 7.0e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.1045e-08+0*(1.1045e-08*(0.02/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.614010248137955+0*(0.0/sqrt(l*w*mult))} lvth0 = -1.01766905880946e-07 wvth0 = -1.93009271144495e-07 pvth0 = 8.83537338381884e-14
+ k1 = 0.825702201038353 lk1 = -9.2805404967024e-08 wk1 = -8.21014511541696e-08 pk1 = 1.80858009105647e-14
+ k2 = -0.0939288954956607 lk2 = 5.54222673537089e-08 wk2 = 2.25615577890959e-08 pk2 = -4.13103838558891e-15
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -35629.1218747767 lvsat = 0.0345810324487428 wvsat = 0.0421601089778771 pvsat = -1.21316102261976e-8
+ ua = -2.01502012646772e-10 lua = 3.8107523195393e-16 wua = -1.6802082660566e-15 pua = 9.22207016602523e-22
+ ub = 2.57984844699042e-18 lub = -1.60283699440755e-25 wub = 4.45694215907796e-24 pub = -2.35603463086626e-30
+ uc = 7.66786672987113e-12 luc = -3.5743851109443e-18 wuc = -1.55955042196236e-18 puc = -3.06700804523122e-25
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0136935482838823 lu0 = -5.17784427064273e-10 wu0 = 2.38986883634779e-09 pu0 = -2.9221952461287e-16
+ a0 = -1.38581975256363 la0 = 1.18012969688866e-06 wa0 = 1.97910647053581e-06 pa0 = -1.04126223230522e-12
+ keta = -0.349400890667415 lketa = 8.89239818704356e-08 wketa = 1.34103041872959e-07 pketa = -3.24414514141805e-14
+ a1 = 0.0
+ a2 = 0.5
+ ags = -1.04896040416374 lags = 1.35686877310111e-06 wags = 1.38455814907852e-06 pags = -9.57728104444705e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {0.00356707220152352+0*(0.009/sqrt(l*w*mult))} lvoff = -4.94492957465713e-08 wvoff = -1.04265205828905e-07 pvoff = 4.71412928422032e-14
+ nfactor = {-3.1691743752861+0*(0.02/sqrt(l*w*mult))} lnfactor = 2.00026493071546e-06 wnfactor = 1.37669490521942e-08 pnfactor = 6.47202997113389e-14
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -5.26977110000001e-05 lcit = 2.34865625406e-11 wcit = 2.8828156726956e-11 pcit = -1.07990275099177e-17
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -1.12297300301366 leta0 = 4.85535502320243e-07 weta0 = 7.15099951647273e-07 peta0 = -2.96967602151934e-13
+ etab = 0.191742400273384 letab = -6.30251871957698e-08 wetab = -1.29733411502351e-07 petab = 4.08751247324909e-14
+ dsub = 0.402842227810149 ldsub = -5.61915155069674e-08 wdsub = -2.53465603885534e-08 pdsub = 1.41593824982339e-14
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 3.15218704400743 lpclm = -8.24127438916613e-07 wpclm = -9.30696290703005e-07 ppclm = 3.72758023840188e-13
+ pdiblc1 = 5.36198413528038 lpdiblc1 = -2.06900528795049e-06 wpdiblc1 = -2.36184826533483e-06 ppdiblc1 = 9.79442875353867e-13
+ pdiblc2 = 0.0380016354791449 lpdiblc2 = -1.48608455845408e-08 wpdiblc2 = -2.24221751084004e-08 ppdiblc2 = 9.88885069851329e-15
+ pdiblcb = -0.025
+ drout = 2.12026187822023 ldrout = -3.12964170720035e-07 wdrout = -8.31829333722917e-07 pdrout = 2.32677444984759e-13
+ pscbe1 = 284930947.001659 lpscbe1 = 66.2950015231527 wpscbe1 = 85.1276251319609 ppscbe1 = -4.90447769468223e-5
+ pscbe2 = 1.8508164228348e-08 lpscbe2 = -1.38570667490259e-15 wpscbe2 = -3.70499341724753e-15 ppscbe2 = 1.36915902245593e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.000150179405180373 lalpha0 = -4.37743113760781e-11 walpha0 = -4.46500989015194e-11 palpha0 = 1.28775076955296e-17
+ alpha1 = 0.0
+ beta0 = 75.0136537213555 lbeta0 = -8.67165998765272e-06 wbeta0 = -1.08988761061372e-05 pbeta0 = 2.62971006543912e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -3.32262249680572e-07 lagidl = 1.31833393900399e-13 wagidl = 2.55972116019088e-13 pagidl = -9.21373027146181e-20
+ bgidl = 2125787493.8811 lbgidl = -58.324672932431 wbgidl = -405.436685619259 pbgidl = 0.000100361626085621
+ cgidl = -8429.85281797858 lcgidl = 0.00351680780080864 wcgidl = 0.00671735716268928 pcgidl = -2.54911044371608e-9
+ egidl = -0.589319140020146 legidl = 4.31455078315809e-07 wegidl = 1.20768668365442e-06 pegidl = -3.50744422241771e-13
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.441061413628573 lkt1 = -7.70838610918801e-08 wkt1 = 4.55079119676261e-09 pkt1 = -2.15980550198351e-15
+ kt2 = -0.019032
+ at = 108698.377171429 lat = -0.0468422498055601 wat = -0.0591602855579143 pat = 2.80774715257861e-8
+ ute = -1.96987764187429 lute = 2.20434986833536e-07 wute = 5.4379743792243e-07 pute = -2.00429950584073e-13
+ ua1 = 5.52e-10
+ ub1 = -1.66079978319999e-19 lub1 = -8.08490602289326e-25 wub1 = 9.81150582022026e-25 pub1 = -4.65654066227653e-31
+ uc1 = 1.2110251937472e-09 luc1 = -5.36203888408582e-16 wuc1 = -7.23647349510653e-16 puc1 = 3.01888973845252e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 1.81e-6
+ sbref = 1.81e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.ends sky130_fd_pr__pfet_g5v0d10v5
