* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
.subckt  sky130_fd_pr__pfet_g5v0d10v5 d g s b
+ 
.param  l = 1 w = 1 ad = 0 as = 0 pd = 0 ps = 0 nrd = 0 nrs = 0 sa = 0 sb = 0 sd = 0 mult = 1 nf = 1.0
msky130_fd_pr__pfet_g5v0d10v5 d g s b sky130_fd_pr__pfet_g5v0d10v5__model l = {l} w = {w} ad = {ad} as = {as} pd = {pd} ps = {ps} nrd = {nrd} nrs = {nrs} sa = {sa} sb = {sb} sd = {sd} nf = {nf}
.model sky130_fd_pr__pfet_g5v0d10v5__model.0 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 2.0e-05 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.042752+0*(0.0/sqrt(l*w*mult))}
+ k1 = 0.59521
+ k2 = 0.0283168
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200000.0
+ ua = 2.7086332e-9
+ ub = -4.1451e-19
+ uc = -3.9972e-11
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0204141
+ a0 = 0.909575
+ keta = -0.0079259
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.120633
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.093204657+0*(0.009/sqrt(l*w*mult))}
+ nfactor = {1.72595+0*(0.02/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.08353125
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0029407877
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 333712830.0
+ pscbe2 = 1.5000958e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 5.0667189e-5
+ alpha1 = 0.0
+ beta0 = 38.266046
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 7.3657e-9
+ bgidl = 1704700000.0
+ cgidl = 700.0
+ egidl = 0.69350825
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.57573
+ kt2 = -0.019032
+ at = 430000.0
+ ute = -1.3864
+ ua1 = 7.0656e-10
+ ub1 = -3.145e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.1 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 2.0e-05 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.042752+0*(0.0/sqrt(l*w*mult))}
+ k1 = 0.59521
+ k2 = 0.0283168
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200000.0
+ ua = 2.7086332e-9
+ ub = -4.1451e-19
+ uc = -3.9972e-11
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0204141
+ a0 = 0.909575
+ keta = -0.0079259
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.120633
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.093204657+0*(0.009/sqrt(l*w*mult))}
+ nfactor = {1.72595+0*(0.02/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.08353125
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0029407877
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 333712830.0
+ pscbe2 = 1.5000958e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 5.0667189e-5
+ alpha1 = 0.0
+ beta0 = 38.266046
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 7.3657e-9
+ bgidl = 1704700000.0
+ cgidl = 700.0
+ egidl = 0.69350825
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.57573
+ kt2 = -0.019032
+ at = 430000.0
+ ute = -1.3864
+ ua1 = 7.0656e-10
+ ub1 = -3.145e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.2 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 2.0e-05 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.04718997701625+0*(0.0/sqrt(l*w*mult))} lvth0 = 3.52087128483047e-8
+ k1 = 0.6042078926875 lk1 = -7.13848266257453e-8
+ k2 = 0.0266281463035 lk2 = 1.33969425444512e-8
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 298327.7912375 lvsat = -0.780084023421662
+ ua = 2.45472545225e-09 lua = 2.01437838631336e-15
+ ub = -1.530400888875e-19 lub = -2.07437284716057e-24
+ uc = -5.164762621625e-11 luc = 9.26286389647505e-17
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.019611959992875 lu0 = 6.36378175722622e-9
+ a0 = 0.9336342833325 la0 = -1.90874444614806e-7
+ keta = -0.004938304614875 lketa = -2.37021029258661e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.0987686124575 lags = 1.73461227890361e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0947862308566375+0*(0.009/sqrt(l*w*mult))} lvoff = 1.25474240995029e-8
+ nfactor = {1.7533173610375+0*(0.02/sqrt(l*w*mult))} lnfactor = -2.17119095627811e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.652860044042275 lpclm = 5.84216401324086e-06 wpclm = 1.6940658945086e-21 ppclm = -9.69352280335579e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00456413311797212 lpdiblc2 = -1.28788189902089e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 563540476.342287 lpscbe1 = -1823.33878139477
+ pscbe2 = -1.55054993344525e-08 lpscbe2 = 2.42023131795166e-13 ppscbe2 = 3.85185988877447e-34
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 7.8323760992625e-05 lalpha0 = -2.1941355218635e-10
+ alpha1 = 0.0
+ beta0 = 39.1457124405462 lbeta0 = -6.97883810440585e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 6.533665354875e-09 lagidl = 6.60095101727241e-15
+ bgidl = 1476950060.5 lbgidl = 1806.85528377295
+ cgidl = 934.0435475 lcgidl = -0.00185678565430899
+ egidl = 1.21251915959209 legidl = -4.11757564630338e-6
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.5852982509125 lkt1 = 7.59097664555738e-8
+ kt2 = -0.019032
+ at = 674555.8396125 lat = -1.94018497634497
+ ute = -1.219521050375 lute = -1.32393498124468e-6
+ ua1 = 1.37964564158e-09 lua1 = -5.33992830290314e-15
+ ub1 = -2.60709319125e-18 lub1 = -4.26748635675217e-24
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.3 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 2.0e-05 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.0234157839175+0*(0.0/sqrt(l*w*mult))} lvth0 = -5.83071945765935e-8
+ k1 = 0.6028041533 lk1 = -6.58632107263166e-8
+ k2 = 0.02903969505375 lk2 = 3.91110347759907e-9
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 84348.6095 lvsat = 0.0616041578387025
+ ua = 3.26941986855725e-09 lua = -1.19022617370328e-15
+ ub = -1.702189719825e-18 lub = 4.01921497188024e-24
+ uc = -5.52637784975e-11 luc = 1.06852792043809e-16
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.02047196271525 lu0 = 2.98095674875055e-9
+ a0 = 0.8170563912675 la0 = 2.67685276712333e-7
+ keta = -0.00501267161 lketa = -2.34095799787069e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.0957090064005 lags = 1.85496203613601e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0637375436500175+0*(0.009/sqrt(l*w*mult))} lvoff = -1.09582742271173e-7
+ nfactor = {2.1038921265675+0*(0.02/sqrt(l*w*mult))} lnfactor = -1.59610668871389e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.0183211905 leta0 = 2.42613905562298e-7
+ etab = -0.12306697823 letab = 2.08739224202596e-7
+ dsub = 0.817977904625 ldsub = -1.01475737773196e-6
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.05151476838812 lpclm = -8.62002833328182e-7
+ pdiblc1 = 0.5839957106185 lpdiblc1 = -7.63083097696423e-7
+ pdiblc2 = -0.00116412829032 lpdiblc2 = 9.65332590061517e-09 ppdiblc2 = -2.52435489670724e-29
+ pdiblcb = 0.1683505 lpdiblcb = -7.605451585025e-07 ppdiblcb = -4.03896783473158e-28
+ drout = 0.1346289 ldrout = 1.6731993487055e-6
+ pscbe1 = -159424727.08145 lpscbe1 = 1020.44846109852 ppscbe1 = -1.73472347597681e-18
+ pscbe2 = 7.64564645311875e-08 lpscbe2 = -1.19709712880149e-13
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 4.43365799732225e-05 lalpha0 = -8.57248057106256e-11
+ alpha1 = -9.667525e-11 lalpha1 = 3.8027257925125e-16
+ beta0 = 70.6002512545225 lbeta0 = -0.000130705423801876
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 9.2096819305e-09 lagidl = -3.9251735630314e-15
+ bgidl = 2628688140.5 lbgidl = -2723.51221259745
+ cgidl = 455.667771125 lcgidl = 2.49078539409564e-5
+ egidl = -1.60756773472605 legidl = 6.97525025293149e-06 wegidl = -3.3881317890172e-21
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.5669667525 lkt1 = 3.8027257925123e-9
+ kt2 = -0.019032
+ at = 210805.618775 lat = -0.116021163929556
+ ute = -1.70701006525 lute = 5.93605496211202e-7
+ ua1 = -4.9057671776e-10 lua1 = 2.01660069867255e-15 wua1 = -5.91645678915759e-31 pua1 = 1.1284745767894e-36
+ ub1 = -3.72032584825e-18 lub1 = 1.11419865720615e-25
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.4 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 2.0e-05 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.0736423575+0*(0.0/sqrt(l*w*mult))} lvth0 = 3.88061365780371e-8
+ k1 = 0.55879817175 lk1 = 1.92225746305162e-8
+ k2 = 0.0262936897075 lk2 = 9.22051854460022e-9
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 179987.995105 lvsat = -0.123315072425493
+ ua = 3.545625841344e-09 lua = -1.72427180311633e-15
+ ub = -3.27932723999998e-20 lub = 7.91428593801762e-25
+ uc = 5.465298373e-13 luc = -1.05671817306874e-18
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.024960961986 lu0 = -5.69854578624093e-9
+ a0 = 1.078927230585 la0 = -2.3864330046225e-7
+ keta = 0.04594012976 lketa = -1.21927076191609e-07 wketa = -1.05879118406788e-22 pketa = 1.0097419586829e-28
+ a1 = 0.0
+ a2 = 0.5
+ ags = -0.268103665696 lags = 8.88929824175545e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.160234189396785+0*(0.009/sqrt(l*w*mult))} lvoff = 7.69940047634308e-8
+ nfactor = {1.017033070615+0*(0.02/sqrt(l*w*mult))} lnfactor = 5.05340730265545e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.4667525e-05 lcit = -9.024682925125e-12
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.278011282483295 leta0 = -2.59498185737863e-7
+ etab = -0.02921139354 letab = 2.72689819265577e-8
+ dsub = 0.0588309099500002 ldsub = 4.53057132207125e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.0480063634240999 lpclm = 1.07828568521179e-6
+ pdiblc1 = -0.00688436326899999 lpdiblc1 = 3.79386479565428e-7
+ pdiblc2 = 0.0059964470822665 lpdiblc2 = -4.19168238515769e-9
+ pdiblcb = -0.411701 lpdiblcb = 3.60987317005e-07 wpdiblcb = -1.6940658945086e-21
+ drout = 1.55012438231795 ldrout = -1.06366824383367e-6
+ pscbe1 = 432633596.7114 lpscbe1 = -124.299268246575
+ pscbe2 = 1.453248063888e-08 lpscbe2 = 2.06195955473267e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -6.3303731508805e-05 lalpha0 = 1.22398274741432e-10 walpha0 = -7.8767761386318e-26 palpha0 = 5.72941588963667e-32
+ alpha1 = 1.933505e-10 lalpha1 = -1.804936585025e-16
+ beta0 = -41.017491252125 lbeta0 = 8.510803942344e-05 wbeta0 = -8.13151629364128e-20 pbeta0 = -1.55096364853693e-25
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 3.753263248e-09 lagidl = 6.62483924167576e-15
+ bgidl = 845577794.0 lbgidl = 724.14055791203
+ cgidl = 438.74318535 lcgidl = 5.76316251598482e-5
+ egidl = 3.1398290592442 legidl = -2.20386518519396e-6
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.498534444 lkt1 = -1.2851148485378e-7
+ kt2 = -0.019032
+ at = 263754.105 lat = -0.218397326788025
+ ute = -1.2068578155 lute = -3.73441379441673e-7
+ ua1 = 6.761640929e-10 lua1 = -2.39298492442614e-16 wua1 = -3.15544362088405e-30
+ ub1 = -3.5285553315e-18 lub1 = -2.59369387268094e-25
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.81e-6
+ sbref = 2.81e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.5 pmos
* DC IV MOS Parameters
+ lmin = 8.0e-07 lmax = 1e-06 wmin = 2.0e-05 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.107061883675+0*(0.0/sqrt(l*w*mult))} lvth0 = 7.0003431360031e-8
+ k1 = 0.5906126265 lk1 = -1.04763779508825e-8
+ k2 = 0.02953277975 lk2 = 6.19681179447626e-9
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 13061.449095 lvsat = 0.032511692907572
+ ua = -8.49051659820001e-10 lua = 2.37818161760777e-15
+ ub = 4.71193868875e-18 lub = -3.63780241559157e-24
+ uc = 6.3107339585e-12 luc = -6.43763154122954e-18
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0179627241575 lu0 = 8.34344217852953e-10
+ a0 = 0.749109306875 la0 = 6.92433804106529e-8
+ keta = -0.15612272205 lketa = 6.66996062872852e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.54854293065 lags = 1.26586143253572e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0958530090713+0*(0.009/sqrt(l*w*mult))} lvoff = 1.68938510236888e-8
+ nfactor = {1.49044010195+0*(0.02/sqrt(l*w*mult))} lnfactor = 6.34128994791644e-8
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -1.3337625e-05 lcit = 1.7118264625625e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -7.5094944625e-05 leta0 = 9.68380229871606e-11
+ etab = 0.00078033929425 letab = -7.28450632878846e-10
+ dsub = 1.5319711835 ldsub = -9.22126678853167e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.04990346593375 lpclm = -7.90495269466486e-7
+ pdiblc1 = 0.18889710180225 lpdiblc1 = 1.96623503014091e-7
+ pdiblc2 = -0.0348197016362825 lpdiblc2 = 3.39103965243514e-08 wpdiblc2 = -2.64697796016969e-23 ppdiblc2 = 2.52435489670724e-29
+ pdiblcb = -0.025
+ drout = 0.3332828474015 ldrout = 7.22594132185131e-8
+ pscbe1 = -69178212.7425001 lpscbe1 = 344.144564937687
+ pscbe2 = 1.840896906885e-08 lpscbe2 = -3.59810173627183e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.00025329086614975 lalpha0 = -1.73144365145817e-10
+ alpha1 = 0.0
+ beta0 = 67.7797653173751 lbeta0 = -1.64547435704711e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 8.97956225e-09 lagidl = 1.74606299181375e-15
+ bgidl = 939140349.999999 lbgidl = 636.799444073251
+ cgidl = 428.889912 lcgidl = 6.68297050984402e-5
+ egidl = 1.87168959037975 legidl = -1.02005065031165e-6
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.6094270675 lkt1 = -2.49926663534123e-8
+ kt2 = -0.019032
+ at = 47404.12 lat = -0.0164335340406
+ ute = -2.0730424275 lute = 4.35146286783388e-7
+ ua1 = -6.64204645000001e-11 lua1 = 4.53907904813073e-16
+ ub1 = -4.5967516375e-18 lub1 = 7.37797205364436e-25
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.41e-6
+ sbref = 2.41e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.6 pmos
* DC IV MOS Parameters
+ lmin = 6e-07 lmax = 8.0e-07 wmin = 2.0e-05 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.946540057525+0*(0.0/sqrt(l*w*mult))} lvth0 = -4.77401307301247e-8
+ k1 = 0.59524275225 lk1 = -1.38725983391364e-8
+ k2 = 0.0329127025 lk2 = 3.7176215577375e-9
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 59860.9299525 lvsat = -0.00181596029880851
+ ua = -2.18776357838e-09 lua = 3.36013350343112e-15
+ ub = 2.580957863135e-18 lub = -2.07471732509884e-24 wub = -2.93873587705572e-39 pub = 4.20389539297445e-45
+ uc = 3.03250253000001e-12 luc = -4.03303239726765e-18
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0061320272125 lu0 = 9.51221958049519e-9
+ a0 = 0.94362221325 la0 = -7.34328089799413e-8
+ keta = 0.0194105553750001 lketa = -6.20549303703394e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = -0.689680622000001 lags = 1.03482931024011e-6
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {0.0153307911677251+0*(0.009/sqrt(l*w*mult))} lvoff = -6.46600223706371e-8
+ nfactor = {1.962272004275+0*(0.02/sqrt(l*w*mult))} lnfactor = -2.82678160035734e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -0.06304090774685 leta0 = 4.62825765424832e-08 weta0 = 1.65436122510606e-23 peta0 = 8.55914082164798e-29
+ etab = -0.00078033929425 letab = 4.16314915178846e-10
+ dsub = 0.1852475514785 ldsub = 6.57018388527629e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.18595238885375 lpclm = 5.76722165327081e-7
+ pdiblc1 = 0.16298765229625 lpdiblc1 = 2.15628213773989e-7
+ pdiblc2 = 0.02744500370811 lpdiblc2 = -1.17610761692872e-8
+ pdiblcb = -0.025
+ drout = -0.7940560006085 ldrout = 8.99168094928088e-7
+ pscbe1 = 433759236.091 lpscbe1 = -24.7625684689289
+ pscbe2 = 1.0404743204925e-08 lpscbe2 = 2.2730379560465e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -0.000128252924521375 lalpha0 = 1.06719913030406e-10 walpha0 = -2.06795153138257e-25 palpha0 = -9.86076131526265e-32
+ alpha1 = 0.0
+ beta0 = 25.56667467665 lbeta0 = 1.45087694799539e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 2.42678867225e-08 lagidl = -9.46799945038737e-15
+ bgidl = 2074319252.5 lbgidl = -195.859956805012
+ cgidl = 1293.58225 lcgidl = -0.00056742644828625
+ egidl = -0.28140889663 legidl = 5.59257855402438e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.7102414755 lkt1 = 4.89552059866275e-8
+ kt2 = -0.019032
+ at = 43672.675 lat = -0.013696500475875
+ ute = -1.6198450625 lute = 1.02723753569062e-7
+ ua1 = 5.5346701e-10 lua1 = -7.82657170049953e-19
+ ub1 = -4.3690170425e-18 lub1 = 5.70752741258962e-25
+ uc1 = -2.898021126e-10 luc1 = 1.32472552602663e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.02e-6
+ sbref = 2.01e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.7 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 6e-07 wmin = 2.0e-05 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.02/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.935589561600001+0*(0.0/sqrt(l*w*mult))} lvth0 = -5.35822750585918e-8
+ k1 = 0.44439056 lk1 = 6.66078004872001e-8
+ k2 = 0.05332399005 lk2 = -7.17190240662526e-9
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 39204.034505 lvsat = 0.00920459670690996
+ ua = 1.2299049456815e-08 lua = -4.36865368491059e-15
+ ub = -1.031258796827e-17 lub = 4.80405384368489e-24
+ uc = -1.256204775e-12 luc = -1.74498560651362e-18
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.03901125958 lu0 = -8.0290152837279e-9
+ a0 = 0.139856216999999 la0 = 3.55380368849415e-7
+ keta = -0.14474227675 lketa = 2.55214263325088e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 1.25
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1246427114985+0*(0.009/sqrt(l*w*mult))} lvoff = 1.00165411693073e-8
+ nfactor = {1.43268543805+0*(0.02/sqrt(l*w*mult))} lnfactor = -1.41079021865146e-10
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 3.167525e-05 lcit = -1.156385425125e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -0.2205430572 leta0 = 1.30310760786486e-07 peta0 = 2.01948391736579e-28
+ etab = 0.016691243015 letab = -8.90486160471758e-9
+ dsub = 0.432939904543 ldsub = -6.64432699689132e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.965059115425 lpclm = 1.61064831167685e-7
+ pdiblc1 = 1.751193186706 lpdiblc1 = -6.31687379861285e-7
+ pdiblc2 = 0.00799763922495 lpdiblc2 = -1.38580998069895e-9
+ pdiblcb = -0.025
+ drout = 0.855521778757 ldrout = 1.91101017476964e-8
+ pscbe1 = 494439169.22 lpscbe1 = -57.1356161929161
+ pscbe2 = 1.54395059094e-08 lpscbe2 = -4.13033120604442e-16
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -3.81232336812e-05 lalpha0 = 5.86352723187186e-11
+ alpha1 = 0.0
+ beta0 = 44.42709312265 lbeta0 = 4.4466419369206e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -2.5414779845e-08 lagidl = 1.70379515767067e-14
+ bgidl = 2109059135.0 lbgidl = -214.393857818175
+ cgidl = -2570.4423 lcgidl = 0.0014940499692615 pcgidl = -1.65436122510606e-24
+ egidl = 1.20727463867 legidl = -2.34962254097789e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.64015525 lkt1 = 1.15638542512501e-8
+ kt2 = -0.019032
+ at = 18000.0
+ ute = -1.665294245 lute = 1.26971119678726e-7
+ ua1 = 5.52e-10
+ ub1 = -8.23768896e-18 lub1 = 2.6347085526048e-24
+ uc1 = -4.1496e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 1.81e-6
+ sbref = 1.81e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.8 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 1.5e-05 wmax = 2.0e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.042752+0*(0.0/sqrt(l*w*mult))}
+ k1 = 0.59521
+ k2 = 0.0283168
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200000.0
+ ua = 2.7086332e-9
+ ub = -4.1451e-19
+ uc = -3.9972e-11
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0204141
+ a0 = 0.909575
+ keta = -0.0079259
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.120633
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.093204657+0*(0.009/sqrt(l*w*mult))}
+ nfactor = {1.72595+0*(0.02/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.08353125
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0029407877
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 333712830.0
+ pscbe2 = 1.5000958e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 5.0667189e-5
+ alpha1 = 0.0
+ beta0 = 38.266046
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 7.3657e-9
+ bgidl = 1704700000.0
+ cgidl = 700.0
+ egidl = 0.69350825
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.57573
+ kt2 = -0.019032
+ at = 430000.0
+ ute = -1.3864
+ ua1 = 7.0656e-10
+ ub1 = -3.145e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.9 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 1.5e-05 wmax = 2.0e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.042752+0*(0.0/sqrt(l*w*mult))}
+ k1 = 0.59521
+ k2 = 0.0283168
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200000.0
+ ua = 2.7086332e-9
+ ub = -4.1451e-19
+ uc = -3.9972e-11
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0204141
+ a0 = 0.909575
+ keta = -0.0079259
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.120633
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.093204657+0*(0.009/sqrt(l*w*mult))}
+ nfactor = {1.72595+0*(0.02/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.08353125
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0029407877
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 333712830.0
+ pscbe2 = 1.5000958e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 5.0667189e-5
+ alpha1 = 0.0
+ beta0 = 38.266046
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 7.3657e-9
+ bgidl = 1704700000.0
+ cgidl = 700.0
+ egidl = 0.69350825
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.57573
+ kt2 = -0.019032
+ at = 430000.0
+ ute = -1.3864
+ ua1 = 7.0656e-10
+ ub1 = -3.145e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.10 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 1.5e-05 wmax = 2.0e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.04718997701625+0*(0.0/sqrt(l*w*mult))} lvth0 = 3.5208712848303e-8
+ k1 = 0.604207892687501 lk1 = -7.13848266257419e-8
+ k2 = 0.0266281463035 lk2 = 1.33969425444513e-8
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 298327.7912375 lvsat = -0.780084023421662
+ ua = 2.45472545225e-09 lua = 2.01437838631335e-15
+ ub = -1.530400888875e-19 lub = -2.07437284716058e-24
+ uc = -5.164762621625e-11 luc = 9.26286389647506e-17
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.019611959992875 lu0 = 6.36378175722624e-9
+ a0 = 0.933634283332501 la0 = -1.90874444614805e-7
+ keta = -0.00493830461487501 lketa = -2.37021029258661e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.0987686124575001 lags = 1.73461227890361e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0947862308566375+0*(0.009/sqrt(l*w*mult))} lvoff = 1.25474240995026e-8
+ nfactor = {1.7533173610375+0*(0.02/sqrt(l*w*mult))} lnfactor = -2.17119095627804e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.652860044042275 lpclm = 5.84216401324086e-06 wpclm = 1.6940658945086e-21 ppclm = -2.58493941422821e-26
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00456413311797213 lpdiblc2 = -1.28788189902089e-08 wpdiblc2 = -5.29395592033938e-23
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 563540476.342287 lpscbe1 = -1823.33878139477
+ pscbe2 = -1.55054993344525e-08 lpscbe2 = 2.42023131795166e-13 ppscbe2 = 1.54074395550979e-33
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 7.8323760992625e-05 lalpha0 = -2.1941355218635e-10
+ alpha1 = 0.0
+ beta0 = 39.1457124405462 lbeta0 = -6.97883810440569e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 6.533665354875e-09 lagidl = 6.6009510172724e-15
+ bgidl = 1476950060.5 lbgidl = 1806.85528377294
+ cgidl = 934.043547499999 lcgidl = -0.00185678565430899
+ egidl = 1.21251915959209 legidl = -4.11757564630337e-6
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.5852982509125 lkt1 = 7.59097664555754e-8
+ kt2 = -0.019032
+ at = 674555.8396125 lat = -1.94018497634497
+ ute = -1.219521050375 lute = -1.32393498124469e-6
+ ua1 = 1.37964564158e-09 lua1 = -5.33992830290314e-15
+ ub1 = -2.60709319125e-18 lub1 = -4.26748635675217e-24
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.11 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 1.5e-05 wmax = 2.0e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.0234157839175+0*(0.0/sqrt(l*w*mult))} lvth0 = -5.83071945765952e-8
+ k1 = 0.6028041533 lk1 = -6.58632107263162e-8
+ k2 = 0.02903969505375 lk2 = 3.91110347759907e-9
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 84348.6095 lvsat = 0.0616041578387025
+ ua = 3.26941986855725e-09 lua = -1.19022617370328e-15
+ ub = -1.702189719825e-18 lub = 4.01921497188023e-24 wub = 1.17549435082229e-38
+ uc = -5.52637784975e-11 luc = 1.06852792043809e-16
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.02047196271525 lu0 = 2.98095674875057e-9
+ a0 = 0.8170563912675 la0 = 2.6768527671233e-7
+ keta = -0.00501267161000001 lketa = -2.34095799787069e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.0957090064005002 lags = 1.85496203613601e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0637375436500175+0*(0.009/sqrt(l*w*mult))} lvoff = -1.09582742271173e-7
+ nfactor = {2.1038921265675+0*(0.02/sqrt(l*w*mult))} lnfactor = -1.59610668871389e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.0183211905 leta0 = 2.42613905562298e-7
+ etab = -0.12306697823 letab = 2.08739224202596e-7
+ dsub = 0.817977904625001 ldsub = -1.01475737773196e-6
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.05151476838812 lpclm = -8.62002833328181e-7
+ pdiblc1 = 0.5839957106185 lpdiblc1 = -7.63083097696422e-7
+ pdiblc2 = -0.00116412829032 lpdiblc2 = 9.65332590061517e-9
+ pdiblcb = 0.1683505 lpdiblcb = -7.605451585025e-07 wpdiblcb = 8.470329472543e-22
+ drout = 0.1346289 ldrout = 1.6731993487055e-6
+ pscbe1 = -159424727.08145 lpscbe1 = 1020.44846109852
+ pscbe2 = 7.64564645311875e-08 lpscbe2 = -1.19709712880149e-13
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 4.43365799732225e-05 lalpha0 = -8.57248057106256e-11
+ alpha1 = -9.667525e-11 lalpha1 = 3.8027257925125e-16
+ beta0 = 70.6002512545226 lbeta0 = -0.000130705423801876
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 9.20968193050001e-09 lagidl = -3.9251735630314e-15
+ bgidl = 2628688140.5 lbgidl = -2723.51221259745
+ cgidl = 455.667771125 lcgidl = 2.49078539409564e-5
+ egidl = -1.60756773472605 legidl = 6.97525025293149e-06 wegidl = 6.7762635780344e-21
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.5669667525 lkt1 = 3.8027257925123e-9
+ kt2 = -0.019032
+ at = 210805.618775 lat = -0.116021163929557
+ ute = -1.70701006525 lute = 5.936054962112e-7
+ ua1 = -4.9057671776e-10 lua1 = 2.01660069867255e-15 wua1 = 7.88860905221012e-31 pua1 = -7.52316384526264e-36
+ ub1 = -3.72032584825e-18 lub1 = 1.11419865720615e-25
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.12 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 1.5e-05 wmax = 2.0e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.05777857133112+0*(0.0/sqrt(l*w*mult))} lvth0 = 8.13342670157949e-09 wvth0 = -3.16171699042938e-07 pvth0 = 6.11319560958029e-13
+ k1 = 0.558798171749999 lk1 = 1.92225746305166e-8
+ k2 = 0.0265473541849851 lk2 = 8.73005700906031e-09 wk2 = -5.05563602405676e-09 pk2 = 9.7750975306942e-15
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 179987.995105 lvsat = -0.123315072425493
+ ua = 3.52426506232237e-09 lua = -1.68297063007411e-15 wua = 4.25728998377455e-16 pua = -8.23149147007805e-22
+ ub = -1.44790655415944e-18 lub = 3.52755719965005e-24 wub = 2.8203782241458e-23 pub = -5.45321539827703e-29
+ uc = 5.465298373e-13 luc = -1.05671817306874e-18
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.021405478018612 lu0 = 1.17600024212353e-09 wu0 = 7.08622389965326e-08 pu0 = -1.37012493410991e-13
+ a0 = 1.09212614597942 la0 = -2.64163469371937e-07 wa0 = -2.63059742570422e-07 pa0 = 5.0862732755862e-13
+ keta = 0.04594012976 lketa = -1.21927076191609e-7
+ a1 = 0.0
+ a2 = 0.5
+ ags = -0.20642138484115 lags = 7.6966682573129e-07 wags = -1.22935290044317e-06 pags = 2.37695997977137e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.160234189396785+0*(0.009/sqrt(l*w*mult))} lvoff = 7.69940047634307e-8
+ nfactor = {1.22149778955495+0*(0.02/sqrt(l*w*mult))} lnfactor = 1.10007173871557e-07 wnfactor = -4.07506486114909e-06 pnfactor = 7.87915828435607e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.4667525e-05 lcit = -9.024682925125e-12
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.27804885270118 leta0 = -2.59570827941995e-07 weta0 = -7.48789695958379e-10 peta0 = 1.4477886210859e-15
+ etab = -0.02921139354 letab = 2.72689819265577e-8
+ dsub = 0.0588309099500002 ldsub = 4.53057132207125e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.0480063634240997 lpclm = 1.07828568521179e-6
+ pdiblc1 = -0.00688436326899966 lpdiblc1 = 3.79386479565428e-7
+ pdiblc2 = 0.0059964470822665 lpdiblc2 = -4.19168238515769e-9
+ pdiblcb = -0.411701 lpdiblcb = 3.60987317005e-7
+ drout = 1.55012438231795 ldrout = -1.06366824383367e-06 wdrout = 1.35525271560688e-20 pdrout = -1.29246970711411e-26
+ pscbe1 = 432633596.7114 lpscbe1 = -124.299268246576
+ pscbe2 = 1.453248063888e-08 lpscbe2 = 2.06195955473393e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -6.3303731508805e-05 lalpha0 = 1.22398274741432e-10 walpha0 = 2.81023808875933e-25 palpha0 = -6.81636260200022e-31
+ alpha1 = 1.933505e-10 lalpha1 = -1.804936585025e-16
+ beta0 = -41.017491252125 lbeta0 = 8.510803942344e-05 wbeta0 = 1.0842021724855e-19 pbeta0 = -2.06795153138257e-25
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -3.22557615674517e-09 lagidl = 2.01184601249476e-14 wagidl = 1.3909110274537e-13 pagidl = -2.68933342613686e-19
+ bgidl = 1034014262.98897 lbgidl = 359.797702939521 wbgidl = -3755.61533215648 pbgidl = 0.00726150102280121
+ cgidl = 69.4523064793175 lcgidl = 0.000771657385910706 wcgidl = 0.00736011714798952 pcgidl = -1.42308233062235e-8
+ egidl = 3.1398290592442 legidl = -2.20386518519396e-06 wegidl = 2.71050543121376e-20 pegidl = -2.58493941422821e-26
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.51247205265303 lkt1 = -1.01563048835103e-07 wkt1 = 2.77782199124005e-07 pkt1 = -5.37093270917252e-13
+ kt2 = -0.019032
+ at = 269329.148461212 lat = -0.229176701195496 wat = -0.1111128796496 pat = 2.14837308366899e-7
+ ute = -1.2068578155 lute = -3.73441379441671e-7
+ ua1 = 6.761640929e-10 lua1 = -2.39298492442614e-16
+ ub1 = -3.5285553315e-18 lub1 = -2.59369387268095e-25
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.81e-6
+ sbref = 2.81e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.13 pmos
* DC IV MOS Parameters
+ lmin = 8.0e-07 lmax = 1e-06 wmin = 1.5e-05 wmax = 2.0e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.18638081451939+0*(0.0/sqrt(l*w*mult))} lvth0 = 1.28184263729049e-07 wvth0 = 1.58085849521469e-06 pvth0 = -1.15956761053249e-12
+ k1 = 0.590612626499999 lk1 = -1.04763779508838e-8
+ k2 = 0.0282644573625742 lk2 = 7.12713260726498e-09 wk2 = 2.52781801202834e-08 pk2 = -1.85416715091292e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 13061.4490949999 lvsat = 0.0325116929075721
+ ua = -7.42247764711837e-10 lua = 2.29984042652645e-15 wua = -2.12864499188723e-15 pua = 1.56137174477427e-21
+ ub = 1.17875050975472e-17 lub = -8.82776575427637e-24 wub = -1.41018911207291e-22 pub = 1.03438076465104e-28
+ uc = 6.31073395850001e-12 luc = -6.43763154122954e-18 puc = 2.35098870164458e-38
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0357401439944398 lu0 = -1.22054821196416e-08 wu0 = -3.54311194982664e-07 pu0 = 2.59889033075759e-13
+ a0 = 0.683114729902902 la0 = 1.17650732592569e-07 wa0 = 1.31529871285211e-06 pa0 = -9.64778182370598e-13
+ keta = -0.15612272205 lketa = 6.66996062872854e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.240131526375752 lags = 3.52807450345755e-07 wags = 6.14676450221588e-06 pags = -4.50868249619786e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0958530090712999+0*(0.009/sqrt(l*w*mult))} lvoff = 1.6893851023689e-8
+ nfactor = {0.468116507250247+0*(0.02/sqrt(l*w*mult))} lnfactor = 8.13292367809406e-07 wnfactor = 2.03753243057455e-05 pnfactor = -1.49454022548858e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -1.3337625e-05 lcit = 1.7118264625625e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -0.000262946034050539 leta0 = 2.3462773633624e-10 weta0 = 3.74394847979329e-09 peta0 = -2.74620492967078e-15
+ etab = 0.00078033929425 letab = -7.28450632878846e-10
+ dsub = 1.5319711835 ldsub = -9.22126678853168e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.04990346593375 lpclm = -7.90495269466485e-7
+ pdiblc1 = 0.18889710180225 lpdiblc1 = 1.96623503014091e-7
+ pdiblc2 = -0.0348197016362825 lpdiblc2 = 3.39103965243514e-08 wpdiblc2 = -1.05879118406788e-22
+ pdiblcb = -0.025
+ drout = 0.333282847401499 ldrout = 7.22594132185127e-8
+ pscbe1 = -69178212.7425003 lpscbe1 = 344.144564937688
+ pscbe2 = 1.840896906885e-08 lpscbe2 = -3.59810173627181e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.00025329086614975 lalpha0 = -1.73144365145817e-10
+ alpha1 = 0.0
+ beta0 = 67.779765317375 lbeta0 = -1.64547435704711e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 4.38737592737259e-08 lagidl = -2.38490049960743e-14 wagidl = -6.9545551372685e-13 pagidl = 5.10120096596213e-19
+ bgidl = -3041994.94483185 lbgidl = 1327.89490500201 wbgidl = 18778.0766607825 pbgidl = -0.0137738131210672
+ cgidl = 2275.34430635342 lcgidl = -0.00128755382543176 wcgidl = -0.0368005857399477 pcgidl = 2.69934136431803e-8
+ egidl = 1.87168959037975 legidl = -1.02005065031165e-6
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.539739024234848 lkt1 = -7.61091945286164e-08 wkt1 = -1.38891099562001e-06 pkt1 = 1.01877315984226e-12
+ kt2 = -0.019032
+ at = 19528.90269394 lat = 0.00401307722948158 wat = 0.555564398248002 pat = -4.07509263936901e-7
+ ute = -2.0730424275 lute = 4.35146286783388e-7
+ ua1 = -6.64204645000009e-11 lua1 = 4.53907904813073e-16
+ ub1 = -4.59675163749999e-18 lub1 = 7.37797205364436e-25
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.41e-6
+ sbref = 2.41e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.14 pmos
* DC IV MOS Parameters
+ lmin = 6e-07 lmax = 8.0e-07 wmin = 1.5e-05 wmax = 2.0e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.946540057524999+0*(0.0/sqrt(l*w*mult))} lvth0 = -4.77401307301255e-8
+ k1 = 0.59524275225 lk1 = -1.38725983391358e-8
+ k2 = 0.0329127025 lk2 = 3.71762155773751e-9
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 59860.9299524999 lvsat = -0.00181596029880848
+ ua = -2.18776357838e-09 lua = 3.36013350343112e-15
+ ub = 2.580957863135e-18 lub = -2.07471732509884e-24 wub = 1.17549435082229e-38 pub = 5.60519385729927e-45
+ uc = 3.03250253000001e-12 luc = -4.03303239726765e-18
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0061320272125 lu0 = 9.5122195804952e-9
+ a0 = 0.94362221325 la0 = -7.34328089799413e-8
+ keta = 0.0194105553750002 lketa = -6.20549303703394e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = -0.689680622000001 lags = 1.03482931024011e-6
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {0.015330791167725+0*(0.009/sqrt(l*w*mult))} lvoff = -6.46600223706372e-8
+ nfactor = {1.962272004275+0*(0.02/sqrt(l*w*mult))} lnfactor = -2.82678160035733e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -0.06304090774685 leta0 = 4.62825765424832e-08 weta0 = 1.45583787809333e-22 peta0 = 6.31088724176809e-29
+ etab = -0.00078033929425 letab = 4.16314915178847e-10
+ dsub = 0.185247551478499 ldsub = 6.57018388527629e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.185952388853748 lpclm = 5.7672216532708e-7
+ pdiblc1 = 0.162987652296249 lpdiblc1 = 2.1562821377399e-7
+ pdiblc2 = 0.02744500370811 lpdiblc2 = -1.17610761692872e-8
+ pdiblcb = -0.025
+ drout = -0.7940560006085 ldrout = 8.99168094928089e-7
+ pscbe1 = 433759236.091 lpscbe1 = -24.7625684689292
+ pscbe2 = 1.0404743204925e-08 lpscbe2 = 2.27303795604647e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -0.000128252924521375 lalpha0 = 1.06719913030406e-10 walpha0 = 8.27180612553028e-25
+ alpha1 = 0.0
+ beta0 = 25.56667467665 lbeta0 = 1.45087694799539e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 2.42678867225e-08 lagidl = -9.46799945038738e-15
+ bgidl = 2074319252.5 lbgidl = -195.859956805012
+ cgidl = 1293.58225 lcgidl = -0.00056742644828625
+ egidl = -0.281408896630001 legidl = 5.59257855402439e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.710241475499998 lkt1 = 4.89552059866273e-8
+ kt2 = -0.019032
+ at = 43672.675 lat = -0.013696500475875
+ ute = -1.6198450625 lute = 1.02723753569063e-7
+ ua1 = 5.5346701e-10 lua1 = -7.8265717005015e-19
+ ub1 = -4.3690170425e-18 lub1 = 5.70752741258963e-25
+ uc1 = -2.898021126e-10 luc1 = 1.32472552602663e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.02e-6
+ sbref = 2.01e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.15 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 6e-07 wmin = 1.5e-05 wmax = 2.0e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.00463718510652+0*(0.0/sqrt(l*w*mult))} lvth0 = -1.67450226797433e-08 wvth0 = 1.3761471698202e-06 pvth0 = -7.34181395834936e-13
+ k1 = 0.44439056 lk1 = 6.66078004872005e-8
+ k2 = 0.0320556650741434 lk2 = 4.17485530961913e-09 wk2 = 4.2388635170876e-07 pk2 = -2.26145488068383e-13
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 38517.959505779 lvsat = 0.00957062114936946 wvsat = 0.0136737532809299 pvsat = -7.29501574414061e-9
+ ua = 1.22625839233658e-08 lua = -4.34919914048778e-15 wua = 7.26772886648546e-16 pua = -3.87736968891471e-22
+ ub = -1.11272049437604e-17 lub = 5.23865607319387e-24 wub = 1.62356470560149e-23 pub = -8.6617988826192e-30
+ uc = -1.25620477500001e-12 luc = -1.74498560651362e-18
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.030518168882094 lu0 = -3.49790893094157e-09 wu0 = 1.69270745804089e-07 pu0 = -9.03067892402107e-14
+ a0 = 0.139856216999998 la0 = 3.55380368849415e-7
+ keta = -0.14474227675 lketa = 2.55214263325087e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 1.25
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1246427114985+0*(0.009/sqrt(l*w*mult))} lvoff = 1.00165411693071e-8
+ nfactor = {6.07637759787291+0*(0.02/sqrt(l*w*mult))} lnfactor = -2.47757406474819e-06 wnfactor = -9.25506700842874e-05 pnfactor = 4.93762452433177e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 3.167525e-05 lcit = -1.156385425125e-11 wcit = 4.13590306276514e-25
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -0.36562850231832 leta0 = 2.07714571184336e-07 weta0 = 2.89161182589885e-06 peta0 = -1.54268936717616e-12
+ etab = 0.016691243015 letab = -8.90486160471757e-9
+ dsub = 0.432939904543 ldsub = -6.64432699689134e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.965059115424999 lpclm = 1.61064831167687e-7
+ pdiblc1 = 1.751193186706 lpdiblc1 = -6.31687379861284e-7
+ pdiblc2 = 0.00799763922494999 lpdiblc2 = -1.38580998069895e-9
+ pdiblcb = -0.025
+ drout = 0.855521778757002 ldrout = 1.91101017476968e-8
+ pscbe1 = 494439169.22 lpscbe1 = -57.1356161929161
+ pscbe2 = 1.54395059094e-08 lpscbe2 = -4.13033120604436e-16
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -3.81232336812e-05 lalpha0 = 5.86352723187186e-11
+ alpha1 = 0.0
+ beta0 = 44.4270931226501 lbeta0 = 4.44664193692074e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -2.82626383323332e-08 lagidl = 1.85572983189914e-14 wagidl = 5.67589758830966e-14 pagidl = -3.02811974285113e-20
+ bgidl = 2173783191.5303 lbgidl = -248.924465597374 wbgidl = -1289.97672461579 pbgidl = 0.000688209032466164
+ cgidl = -9810.73415970548 lcgidl = 0.00535678187787367 wcgidl = 0.144301956322425 pcgidl = -7.69858152077955e-8
+ egidl = 1.20727463867 legidl = -2.34962254097789e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.5107071369394 lkt1 = -5.74973613071451e-08 wkt1 = -2.57995344923165e-06 pkt1 = 1.37641806493235e-12
+ kt2 = -0.019032
+ at = 18000.0
+ ute = -1.665294245 lute = 1.26971119678726e-7
+ ua1 = 5.52e-10
+ ub1 = -8.23768896e-18 lub1 = 2.6347085526048e-24
+ uc1 = -4.1496e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 1.81e-6
+ sbref = 1.81e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.16 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 1.0e-05 wmax = 1.5e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.042752+0*(0.0/sqrt(l*w*mult))}
+ k1 = 0.59521
+ k2 = 0.0283168
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200000.0
+ ua = 2.7086332e-9
+ ub = -4.1451e-19
+ uc = -3.9972e-11
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0204141
+ a0 = 0.909575
+ keta = -0.0079259
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.120633
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.093204657+0*(0.009/sqrt(l*w*mult))}
+ nfactor = {1.72595+0*(0.02/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.08353125
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0029407877
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 333712830.0
+ pscbe2 = 1.5000958e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 5.0667189e-5
+ alpha1 = 0.0
+ beta0 = 38.266046
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 7.3657e-9
+ bgidl = 1704700000.0
+ cgidl = 700.0
+ egidl = 0.69350825
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.57573
+ kt2 = -0.019032
+ at = 430000.0
+ ute = -1.3864
+ ua1 = 7.0656e-10
+ ub1 = -3.145e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.17 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 1.0e-05 wmax = 1.5e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.042752+0*(0.0/sqrt(l*w*mult))}
+ k1 = 0.59521
+ k2 = 0.0283168
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200000.0
+ ua = 2.7086332e-9
+ ub = -4.1451e-19
+ uc = -3.9972e-11
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0204141
+ a0 = 0.909575
+ keta = -0.0079259
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.120633
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.093204657+0*(0.009/sqrt(l*w*mult))}
+ nfactor = {1.72595+0*(0.02/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.08353125
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0029407877
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 333712830.0
+ pscbe2 = 1.5000958e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 5.0667189e-5
+ alpha1 = 0.0
+ beta0 = 38.266046
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 7.3657e-9
+ bgidl = 1704700000.0
+ cgidl = 700.0
+ egidl = 0.69350825
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.57573
+ kt2 = -0.019032
+ at = 430000.0
+ ute = -1.3864
+ ua1 = 7.0656e-10
+ ub1 = -3.145e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.18 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 1.0e-05 wmax = 1.5e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.04718997701625+0*(0.0/sqrt(l*w*mult))} lvth0 = 3.52087128483064e-8
+ k1 = 0.6042078926875 lk1 = -7.13848266257436e-8
+ k2 = 0.0266281463035 lk2 = 1.33969425444513e-8
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 298327.7912375 lvsat = -0.780084023421662
+ ua = 2.45472545225e-09 lua = 2.01437838631337e-15
+ ub = -1.53040088887501e-19 lub = -2.07437284716057e-24
+ uc = -5.164762621625e-11 luc = 9.26286389647506e-17
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.019611959992875 lu0 = 6.36378175722624e-9
+ a0 = 0.9336342833325 la0 = -1.90874444614805e-7
+ keta = -0.004938304614875 lketa = -2.37021029258661e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.0987686124575 lags = 1.73461227890361e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0947862308566376+0*(0.009/sqrt(l*w*mult))} lvoff = 1.25474240995026e-8
+ nfactor = {1.7533173610375+0*(0.02/sqrt(l*w*mult))} lnfactor = -2.17119095627811e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.652860044042275 lpclm = 5.84216401324086e-06 wpclm = -1.6940658945086e-21
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00456413311797213 lpdiblc2 = -1.28788189902089e-08 wpdiblc2 = -2.64697796016969e-23
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 563540476.342288 lpscbe1 = -1823.33878139477
+ pscbe2 = -1.55054993344525e-08 lpscbe2 = 2.42023131795165e-13
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 7.8323760992625e-05 lalpha0 = -2.1941355218635e-10
+ alpha1 = 0.0
+ beta0 = 39.1457124405463 lbeta0 = -6.9788381044058e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 6.533665354875e-09 lagidl = 6.60095101727242e-15
+ bgidl = 1476950060.5 lbgidl = 1806.85528377294
+ cgidl = 934.0435475 lcgidl = -0.00185678565430899
+ egidl = 1.21251915959209 legidl = -4.11757564630338e-06 wegidl = 6.7762635780344e-21
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.5852982509125 lkt1 = 7.59097664555721e-8
+ kt2 = -0.019032
+ at = 674555.8396125 lat = -1.94018497634497
+ ute = -1.219521050375 lute = -1.32393498124468e-6
+ ua1 = 1.37964564158e-09 lua1 = -5.33992830290314e-15
+ ub1 = -2.60709319125e-18 lub1 = -4.26748635675218e-24
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.19 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 1.0e-05 wmax = 1.5e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.0234157839175+0*(0.0/sqrt(l*w*mult))} lvth0 = -5.83071945765935e-8
+ k1 = 0.602804153300001 lk1 = -6.58632107263162e-8
+ k2 = 0.02903969505375 lk2 = 3.91110347759907e-9
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 84348.6095 lvsat = 0.0616041578387023
+ ua = 3.26941986855725e-09 lua = -1.19022617370329e-15
+ ub = -1.702189719825e-18 lub = 4.01921497188024e-24
+ uc = -5.52637784975e-11 luc = 1.06852792043809e-16
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.02047196271525 lu0 = 2.98095674875057e-9
+ a0 = 0.817056391267501 la0 = 2.67685276712333e-7
+ keta = -0.00501267161000001 lketa = -2.3409579978707e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.0957090064005002 lags = 1.85496203613602e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0637375436500175+0*(0.009/sqrt(l*w*mult))} lvoff = -1.09582742271173e-7
+ nfactor = {2.1038921265675+0*(0.02/sqrt(l*w*mult))} lnfactor = -1.59610668871389e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.0183211905000001 leta0 = 2.42613905562298e-7
+ etab = -0.12306697823 letab = 2.08739224202596e-7
+ dsub = 0.817977904625 ldsub = -1.01475737773196e-6
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.05151476838813 lpclm = -8.62002833328181e-7
+ pdiblc1 = 0.5839957106185 lpdiblc1 = -7.63083097696423e-7
+ pdiblc2 = -0.00116412829032 lpdiblc2 = 9.65332590061517e-9
+ pdiblcb = 0.1683505 lpdiblcb = -7.605451585025e-7
+ drout = 0.1346289 ldrout = 1.6731993487055e-6
+ pscbe1 = -159424727.08145 lpscbe1 = 1020.44846109852
+ pscbe2 = 7.64564645311875e-08 lpscbe2 = -1.19709712880149e-13 wpscbe2 = -4.03896783473158e-28
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 4.43365799732225e-05 lalpha0 = -8.57248057106256e-11
+ alpha1 = -9.667525e-11 lalpha1 = 3.8027257925125e-16
+ beta0 = 70.6002512545225 lbeta0 = -0.000130705423801876
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 9.2096819305e-09 lagidl = -3.92517356303139e-15
+ bgidl = 2628688140.5 lbgidl = -2723.51221259745 wbgidl = 1.45519152283669e-11
+ cgidl = 455.667771125 lcgidl = 2.49078539409572e-5
+ egidl = -1.60756773472605 legidl = 6.97525025293149e-06 pegidl = 6.46234853557053e-27
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.5669667525 lkt1 = 3.8027257925123e-9
+ kt2 = -0.019032
+ at = 210805.618775 lat = -0.116021163929556
+ ute = -1.70701006525 lute = 5.93605496211204e-7
+ ua1 = -4.9057671776e-10 lua1 = 2.01660069867255e-15 wua1 = 1.97215226305253e-31
+ ub1 = -3.72032584825e-18 lub1 = 1.11419865720615e-25
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.20 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 1.0e-05 wmax = 1.5e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.06224838969551+0*(0.0/sqrt(l*w*mult))} lvth0 = 1.67758428582153e-08 wvth0 = -2.49435496116366e-07 pvth0 = 4.8228477891847e-13
+ k1 = 0.55879817175 lk1 = 1.92225746305162e-8
+ k2 = 0.025239090002393 lk2 = 1.1259592347423e-08 wk2 = 1.44772793773012e-08 pk2 = -2.79918920624088e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 179987.995105 lvsat = -0.123315072425493
+ ua = 3.54415255031149e-09 lua = -1.72142318753852e-15 wua = 1.28800728379694e-16 pua = -2.49036852325771e-22
+ ub = 9.35409276446867e-19 lub = -1.0805958754064e-24 wub = -7.38009073572134e-24 pub = 1.42694423379709e-29
+ uc = 5.465298373e-13 luc = -1.05671817306874e-18
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0267773782600795 lu0 = -9.21059573425507e-09 wu0 = -9.34241260007474e-09 pu0 = 1.80636014743078e-14
+ a0 = 1.05135783151165 la0 = -1.8533772950694e-07 wa0 = 3.45627744368989e-07 pa0 = -6.68272971876164e-13
+ keta = 0.04594012976 lketa = -1.21927076191609e-7
+ a1 = 0.0
+ a2 = 0.5
+ ags = -0.329164850946096 lags = 1.00699193116253e-06 wags = 6.03256882350905e-07 pags = -1.16640019830988e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.160234189396785+0*(0.009/sqrt(l*w*mult))} lvoff = 7.69940047634308e-8
+ nfactor = {0.924773444211325+0*(0.02/sqrt(l*w*mult))} lnfactor = 6.83725179215184e-07 wnfactor = 3.55150084915435e-07 pnfactor = -6.86684464934426e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.4667525e-05 lcit = -9.024682925125e-12
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.277998700702905 leta0 = -2.5947385880257e-7
+ etab = -0.02921139354 letab = 2.72689819265577e-8
+ dsub = 0.05883090995 ldsub = 4.53057132207125e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.0480295386332323 lpclm = 1.07824087582905e-06 wpclm = -3.46015281483842e-10 ppclm = 6.69022276831838e-16
+ pdiblc1 = -0.0068843632690001 lpdiblc1 = 3.79386479565428e-7
+ pdiblc2 = 0.0059964470822665 lpdiblc2 = -4.19168238515769e-9
+ pdiblcb = -0.411701 lpdiblcb = 3.60987317005e-7
+ drout = 1.55012438231795 ldrout = -1.06366824383367e-6
+ pscbe1 = 432633596.7114 lpscbe1 = -124.299268246575
+ pscbe2 = 1.453248063888e-08 lpscbe2 = 2.06195955473393e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -6.3303731508805e-05 lalpha0 = 1.22398274741432e-10 walpha0 = -1.22420957298533e-25 palpha0 = 2.19635759196905e-31
+ alpha1 = 1.933505e-10 lalpha1 = -1.804936585025e-16
+ beta0 = -41.017491252125 lbeta0 = 8.510803942344e-05 wbeta0 = -5.42101086242752e-20 pbeta0 = -1.55096364853693e-25
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 6.09038636600001e-09 lagidl = 2.10600000740717e-15
+ bgidl = 782472856.0 lbgidl = 846.15427105972
+ cgidl = 562.41392775 lcgidl = -0.000181486373624264 wcgidl = 3.46944695195361e-18
+ egidl = 3.1398290592442 legidl = -2.20386518519396e-6
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.473101931617213 lkt1 = -1.77685374708461e-07 wkt1 = -3.10029692209895e-07 pkt1 = 5.99443960036286e-13
+ kt2 = -0.019032
+ at = 258549.864884909 lat = -0.208334902504296 wat = 0.0498262005337331 pat = -9.6339207862974e-8
+ ute = -0.935985971158463 lute = -8.97173444835255e-07 wute = -4.04422660998794e-06 pute = 7.81953237154475e-12
+ ua1 = 9.21969631043744e-10 lua1 = -7.14564729471234e-16 wua1 = -3.66997648153458e-15 pua1 = 7.09591787692952e-21
+ ub1 = -3.12901472605441e-18 lub1 = -1.03188314560018e-24 wub1 = -5.96530345278855e-24 pub1 = 1.15339440524838e-29
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.81e-6
+ sbref = 2.81e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.21 pmos
* DC IV MOS Parameters
+ lmin = 8.0e-07 lmax = 1e-06 wmin = 1.0e-05 wmax = 1.5e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.16403172269745+0*(0.0/sqrt(l*w*mult))} lvth0 = 1.11791093132196e-07 wvth0 = 1.24717748058181e-06 pvth0 = -9.14810917894174e-13
+ k1 = 0.5906126265 lk1 = -1.04763779508812e-8
+ k2 = 0.0348057782755347 lk2 = 2.32904101100387e-09 wk2 = -7.23863968865061e-08 pk2 = 5.30957840482369e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 13061.4490949999 lvsat = 0.0325116929075719
+ ua = -8.41685204657454e-10 lua = 2.37277828591377e-15 wua = -6.44003641898444e-16 pua = 4.72379891350746e-22
+ ub = -1.29074055484326e-19 lub = -8.68953626319692e-26 wub = 3.69004536786066e-23 pub = -2.70666672755263e-29
+ uc = 6.3107339585e-12 luc = -6.43763154122954e-18 puc = 1.17549435082229e-38
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.00888064278710235 lu0 = 7.49609631344651e-09 wu0 = 4.67120630003745e-08 pu0 = -3.42635317710894e-14
+ a0 = 0.886956302241733 la0 = -3.18680799258218e-08 wa0 = -1.72813872184495e-06 pa0 = 1.26759839316688e-12
+ keta = -0.15612272205 lketa = 6.66996062872853e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.853848856900482 lags = -9.73572801807883e-08 wags = -3.01628441175452e-06 pags = 2.21245969744399e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0958530090712998+0*(0.009/sqrt(l*w*mult))} lvoff = 1.68938510236889e-8
+ nfactor = {1.95173823396838+0*(0.02/sqrt(l*w*mult))} lnfactor = -2.74951586846973e-07 wnfactor = -1.77575042457722e-06 pnfactor = 1.3025218151795e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -1.3337625e-05 lcit = 1.7118264625625e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -1.2186042675e-05 leta0 = 5.06940288623259e-11
+ etab = 0.00078033929425 letab = -7.28450632878846e-10
+ dsub = 1.5319711835 ldsub = -9.22126678853167e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.04978758988809 lpclm = -7.90410273807609e-07 wpclm = 1.73007640741243e-09 ppclm = -1.26901969522439e-15
+ pdiblc1 = 0.18889710180225 lpdiblc1 = 1.96623503014091e-7
+ pdiblc2 = -0.0348197016362825 lpdiblc2 = 3.39103965243514e-08 wpdiblc2 = -7.94093388050907e-23 ppdiblc2 = -2.52435489670724e-29
+ pdiblcb = -0.025
+ drout = 0.333282847401501 ldrout = 7.22594132185127e-8
+ pscbe1 = -69178212.7424994 lpscbe1 = 344.144564937687
+ pscbe2 = 1.840896906885e-08 lpscbe2 = -3.59810173627181e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.00025329086614975 lalpha0 = -1.73144365145817e-10
+ alpha1 = 0.0
+ beta0 = 67.7797653173751 lbeta0 = -1.64547435704712e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -2.70605334000001e-09 lagidl = 1.03175204551567e-14
+ bgidl = 1254665040 lbgidl = 405.360506334804
+ cgidl = -189.4638 lcgidl = 0.000520395244619
+ egidl = 1.87168959037975 legidl = -1.02005065031165e-6
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.736589629413936 lkt1 = 6.82817086232697e-08 wkt1 = 1.55014846104944e-06 pkt1 = -1.13704164692207e-12
+ kt2 = -0.019032
+ at = 73425.320575454 lat = -0.0355202147686983 wat = -0.249131002668662 pat = 1.82738836112477e-7
+ ute = -3.42740164920768 lute = 1.42857554770208e-06 wute = 2.02211330499397e-05 pute = -1.4832302197796e-11
+ ua1 = -1.29544815521872e-09 lua1 = 1.3554058610937e-15 wua1 = 1.83498824076729e-14 pua1 = -1.34597304954401e-20
+ ub1 = -6.59445466472797e-18 lub1 = 2.20312236435129e-24 wub1 = 2.98265172639425e-23 pub1 = -2.18778995456882e-29
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.41e-6
+ sbref = 2.41e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.22 pmos
* DC IV MOS Parameters
+ lmin = 6e-07 lmax = 8.0e-07 wmin = 1.0e-05 wmax = 1.5e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.946540057524999+0*(0.0/sqrt(l*w*mult))} lvth0 = -4.77401307301255e-8
+ k1 = 0.59524275225 lk1 = -1.38725983391362e-8
+ k2 = 0.0329127025 lk2 = 3.71762155773751e-9
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 59860.9299524999 lvsat = -0.00181596029880848
+ ua = -2.18776357838e-09 lua = 3.36013350343113e-15
+ ub = 2.580957863135e-18 lub = -2.07471732509884e-24 wub = 5.87747175411144e-39
+ uc = 3.03250253e-12 luc = -4.03303239726765e-18
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0061320272125 lu0 = 9.5122195804952e-9
+ a0 = 0.94362221325 la0 = -7.34328089799405e-8
+ keta = 0.019410555375 lketa = -6.20549303703394e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = -0.689680622000003 lags = 1.03482931024011e-6
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {0.015330791167725+0*(0.009/sqrt(l*w*mult))} lvoff = -6.46600223706372e-8
+ nfactor = {1.962272004275+0*(0.02/sqrt(l*w*mult))} lnfactor = -2.82678160035735e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -0.06304090774685 leta0 = 4.62825765424832e-08 weta0 = 2.15066959263787e-23 peta0 = -9.03245736478059e-29
+ etab = -0.00078033929425 letab = 4.16314915178846e-10
+ dsub = 0.1852475514785 ldsub = 6.57018388527629e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.185952388853748 lpclm = 5.76722165327081e-7
+ pdiblc1 = 0.162987652296249 lpdiblc1 = 2.15628213773989e-7
+ pdiblc2 = 0.02744500370811 lpdiblc2 = -1.17610761692872e-8
+ pdiblcb = -0.025
+ drout = -0.794056000608499 ldrout = 8.99168094928088e-7
+ pscbe1 = 433759236.091001 lpscbe1 = -24.7625684689292
+ pscbe2 = 1.0404743204925e-08 lpscbe2 = 2.2730379560465e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -0.000128252924521375 lalpha0 = 1.06719913030406e-10
+ alpha1 = 0.0
+ beta0 = 25.56667467665 lbeta0 = 1.45087694799539e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 2.42678867225e-08 lagidl = -9.46799945038736e-15
+ bgidl = 2074319252.5 lbgidl = -195.859956805012
+ cgidl = 1293.58225 lcgidl = -0.00056742644828625 wcgidl = 6.93889390390723e-18
+ egidl = -0.281408896630001 legidl = 5.59257855402439e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.710241475500001 lkt1 = 4.89552059866273e-8
+ kt2 = -0.019032
+ at = 43672.675 lat = -0.013696500475875
+ ute = -1.6198450625 lute = 1.02723753569065e-7
+ ua1 = 5.53467010000001e-10 lua1 = -7.8265717005015e-19
+ ub1 = -4.3690170425e-18 lub1 = 5.70752741258963e-25
+ uc1 = -2.898021126e-10 luc1 = 1.32472552602663e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.02e-6
+ sbref = 2.01e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.23 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 6e-07 wmin = 1.0e-05 wmax = 1.5e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.787452670736009+0*(0.0/sqrt(l*w*mult))} lvth0 = -1.32614047018986e-07 wvth0 = -1.86650580664448e-06 pvth0 = 9.95790180373863e-13
+ k1 = 0.44439056 lk1 = 6.66078004872005e-8
+ k2 = 0.0759009987443776 lk2 = -1.92168494301193e-08 wk2 = -2.30742281193306e-07 pk2 = 1.23102160728035e-13
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 66865.3526522378 lvsat = -0.00555285483123213 wvsat = -0.409564335437322 pvsat = 2.18504620777488e-7
+ ua = 1.23160569297125e-08 lua = -4.37772725673876e-15 wua = -7.16008081475152e-17 pua = 3.81993891507233e-23
+ ub = -9.88792430185371e-18 lub = 4.57749365433347e-24 wub = -2.26731607559194e-24 pub = 1.20962446290868e-30
+ uc = -1.25620477500001e-12 luc = -1.74498560651362e-18
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0404374581978919 lu0 = -8.7898993773663e-09 wu0 = 2.11717290877646e-08 pu0 = -1.12952233269679e-14
+ a0 = 0.139856217 la0 = 3.55380368849415e-7
+ keta = -0.14474227675 lketa = 2.55214263325087e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 1.25
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1246427114985+0*(0.009/sqrt(l*w*mult))} lvoff = 1.00165411693074e-8
+ nfactor = {-1.91902594018554+0*(0.02/sqrt(l*w*mult))} lnfactor = 1.78801369982369e-06 wnfactor = 2.68239508727617e-05 pnfactor = -1.43107119103728e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 3.167525e-05 lcit = -1.156385425125e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -0.213308500353006 leta0 = 1.26451088535831e-07 weta0 = 6.17412354635907e-07 peta0 = -3.29392578260029e-13
+ etab = -0.0131441628388898 letab = 7.01247659536189e-09 wetab = 4.45454722573351e-07 petab = -2.37652321766495e-13
+ dsub = 0.432939904543 ldsub = -6.64432699689134e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.0446756318071877 lpclm = 6.52094021595207e-07 wpclm = 1.37416990861083e-05 ppclm = -7.33126517093423e-12
+ pdiblc1 = 1.751193186706 lpdiblc1 = -6.31687379861284e-7
+ pdiblc2 = 0.00799763922494999 lpdiblc2 = -1.38580998069895e-9
+ pdiblcb = -0.025
+ drout = 0.855521778757 ldrout = 1.9110101747696e-8
+ pscbe1 = 494439169.219999 lpscbe1 = -57.1356161929161
+ pscbe2 = 1.54395059094e-08 lpscbe2 = -4.13033120604461e-16
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -3.81232336812002e-05 lalpha0 = 5.86352723187185e-11
+ alpha1 = 0.0
+ beta0 = 44.42709312265 lbeta0 = 4.44664193692068e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -7.75660765807781e-08 lagidl = 4.48609291417281e-14 wagidl = 7.92879326128309e-13 pagidl = -4.23005084886083e-19
+ bgidl = 1550995755.63246 lbgidl = 83.3357453913031 wbgidl = 8008.49254503788 pbgidl = -0.00427257081524043
+ cgidl = -595.191674176333 lcgidl = 0.000440243884131445 wcgidl = 0.00671016550322596 pcgidl = -3.57990684679856e-9
+ egidl = 1.20727463867 legidl = -2.34962254097788e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.68350575 lkt1 = 3.46915627537496e-8
+ kt2 = -0.019032
+ at = 18000.0
+ ute = -1.665294245 lute = 1.26971119678723e-7
+ ua1 = 5.52e-10
+ ub1 = -8.23768896e-18 lub1 = 2.6347085526048e-24
+ uc1 = -4.1496e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 1.81e-6
+ sbref = 1.81e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.24 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 7e-06 wmax = 1.0e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.042752+0*(0.0/sqrt(l*w*mult))}
+ k1 = 0.59521
+ k2 = 0.0283168
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200000.0
+ ua = 2.7086332e-9
+ ub = -4.1451e-19
+ uc = -3.9972e-11
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0204141
+ a0 = 0.909575
+ keta = -0.0079259
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.120633
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.093204657+0*(0.009/sqrt(l*w*mult))}
+ nfactor = {1.72595+0*(0.02/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.08353125
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0029407877
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 333712830.0
+ pscbe2 = 1.5000958e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 5.0667189e-5
+ alpha1 = 0.0
+ beta0 = 38.266046
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 7.3657e-9
+ bgidl = 1704700000.0
+ cgidl = 700.0
+ egidl = 0.69350825
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.57573
+ kt2 = -0.019032
+ at = 430000.0
+ ute = -1.3864
+ ua1 = 7.0656e-10
+ ub1 = -3.145e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.25 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 7e-06 wmax = 1.0e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.042752+0*(0.0/sqrt(l*w*mult))}
+ k1 = 0.59521
+ k2 = 0.0283168
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200000.0
+ ua = 2.7086332e-9
+ ub = -4.1451e-19
+ uc = -3.9972e-11
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0204141
+ a0 = 0.909575
+ keta = -0.0079259
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.120633
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.093204657+0*(0.009/sqrt(l*w*mult))}
+ nfactor = {1.72595+0*(0.02/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.08353125
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0029407877
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 333712830.0
+ pscbe2 = 1.5000958e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 5.0667189e-5
+ alpha1 = 0.0
+ beta0 = 38.266046
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 7.3657e-9
+ bgidl = 1704700000.0
+ cgidl = 700.0
+ egidl = 0.69350825
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.57573
+ kt2 = -0.019032
+ at = 430000.0
+ ute = -1.3864
+ ua1 = 7.0656e-10
+ ub1 = -3.145e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.26 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 7e-06 wmax = 1.0e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.04718997701625+0*(0.0/sqrt(l*w*mult))} lvth0 = 3.5208712848303e-8
+ k1 = 0.6042078926875 lk1 = -7.13848266257453e-8
+ k2 = 0.0266281463035 lk2 = 1.33969425444513e-8
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 298327.7912375 lvsat = -0.780084023421662
+ ua = 2.45472545225e-09 lua = 2.01437838631337e-15
+ ub = -1.530400888875e-19 lub = -2.07437284716057e-24
+ uc = -5.164762621625e-11 luc = 9.26286389647506e-17
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.019611959992875 lu0 = 6.36378175722624e-9
+ a0 = 0.9336342833325 la0 = -1.90874444614808e-7
+ keta = -0.00493830461487501 lketa = -2.37021029258661e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.0987686124575 lags = 1.73461227890361e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0947862308566375+0*(0.009/sqrt(l*w*mult))} lvoff = 1.25474240995026e-8
+ nfactor = {1.7533173610375+0*(0.02/sqrt(l*w*mult))} lnfactor = -2.17119095627811e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.652860044042275 lpclm = 5.84216401324086e-06 wpclm = -8.470329472543e-22 ppclm = 9.69352280335579e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00456413311797213 lpdiblc2 = -1.28788189902089e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 563540476.342288 lpscbe1 = -1823.33878139477
+ pscbe2 = -1.55054993344525e-08 lpscbe2 = 2.42023131795165e-13 ppscbe2 = 3.85185988877447e-34
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 7.8323760992625e-05 lalpha0 = -2.1941355218635e-10
+ alpha1 = 0.0
+ beta0 = 39.1457124405463 lbeta0 = -6.9788381044059e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 6.533665354875e-09 lagidl = 6.60095101727242e-15
+ bgidl = 1476950060.5 lbgidl = 1806.85528377294
+ cgidl = 934.043547499999 lcgidl = -0.00185678565430899
+ egidl = 1.21251915959209 legidl = -4.11757564630338e-6
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.5852982509125 lkt1 = 7.59097664555721e-8
+ kt2 = -0.019032
+ at = 674555.8396125 lat = -1.94018497634497
+ ute = -1.219521050375 lute = -1.32393498124468e-6
+ ua1 = 1.37964564158e-09 lua1 = -5.33992830290314e-15
+ ub1 = -2.60709319125e-18 lub1 = -4.26748635675218e-24
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.27 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 7e-06 wmax = 1.0e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.0234157839175+0*(0.0/sqrt(l*w*mult))} lvth0 = -5.83071945765952e-8
+ k1 = 0.6028041533 lk1 = -6.5863210726317e-8
+ k2 = 0.02903969505375 lk2 = 3.91110347759912e-9
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 84348.6095 lvsat = 0.0616041578387025
+ ua = 3.26941986855725e-09 lua = -1.19022617370329e-15
+ ub = -1.702189719825e-18 lub = 4.01921497188024e-24
+ uc = -5.52637784975e-11 luc = 1.06852792043809e-16
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.02047196271525 lu0 = 2.98095674875057e-9
+ a0 = 0.8170563912675 la0 = 2.67685276712333e-7
+ keta = -0.00501267161000001 lketa = -2.34095799787069e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.0957090064005001 lags = 1.85496203613601e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0637375436500176+0*(0.009/sqrt(l*w*mult))} lvoff = -1.09582742271173e-7
+ nfactor = {2.1038921265675+0*(0.02/sqrt(l*w*mult))} lnfactor = -1.5961066887139e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.0183211905000001 leta0 = 2.42613905562297e-7
+ etab = -0.12306697823 letab = 2.08739224202596e-7
+ dsub = 0.817977904625 ldsub = -1.01475737773196e-06 wdsub = -3.3881317890172e-21
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.05151476838812 lpclm = -8.62002833328181e-7
+ pdiblc1 = 0.5839957106185 lpdiblc1 = -7.63083097696422e-7
+ pdiblc2 = -0.00116412829032 lpdiblc2 = 9.65332590061517e-09 ppdiblc2 = 1.26217744835362e-29
+ pdiblcb = 0.1683505 lpdiblcb = -7.60545158502501e-07 ppdiblcb = 4.03896783473158e-28
+ drout = 0.1346289 ldrout = 1.6731993487055e-6
+ pscbe1 = -159424727.08145 lpscbe1 = 1020.44846109852
+ pscbe2 = 7.64564645311875e-08 lpscbe2 = -1.19709712880149e-13
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 4.43365799732225e-05 lalpha0 = -8.57248057106256e-11
+ alpha1 = -9.667525e-11 lalpha1 = 3.8027257925125e-16
+ beta0 = 70.6002512545225 lbeta0 = -0.000130705423801876
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 9.2096819305e-09 lagidl = -3.9251735630314e-15
+ bgidl = 2628688140.5 lbgidl = -2723.51221259746
+ cgidl = 455.667771125 lcgidl = 2.49078539409564e-5
+ egidl = -1.60756773472605 legidl = 6.97525025293149e-06 wegidl = 8.470329472543e-22 pegidl = -4.8467614016779e-27
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.5669667525 lkt1 = 3.80272579251145e-9
+ kt2 = -0.019032
+ at = 210805.618775 lat = -0.116021163929557
+ ute = -1.70701006525 lute = 5.93605496211204e-7
+ ua1 = -4.9057671776e-10 lua1 = 2.01660069867255e-15 wua1 = -3.94430452610506e-31 pua1 = 1.50463276905253e-36
+ ub1 = -3.72032584825e-18 lub1 = 1.11419865720621e-25
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.28 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 7e-06 wmax = 1.0e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.08736674801+0*(0.0/sqrt(l*w*mult))} lvth0 = 6.53423142510758e-8
+ k1 = 0.55879817175 lk1 = 1.92225746305162e-8
+ k2 = 0.0266969638675 lk2 = 8.4407859398694e-9
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 179987.995105 lvsat = -0.123315072425493
+ ua = 3.557122888924e-09 lua = -1.7465014020975e-15
+ ub = 1.9222810785e-19 lub = 3.56348629981485e-25
+ uc = 5.465298373e-13 luc = -1.05671817306874e-18
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.025836589676 lu0 = -7.39157630299439e-9
+ a0 = 1.08616282784 la0 = -2.5263336393278e-7
+ keta = 0.04594012976 lketa = -1.21927076191609e-07 pketa = 2.01948391736579e-28
+ a1 = 0.0
+ a2 = 0.5
+ ags = -0.268416389871 lags = 8.89534477931528e-07 pags = 1.61558713389263e-27
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.160234189396785+0*(0.009/sqrt(l*w*mult))} lvoff = 7.69940047634309e-8
+ nfactor = {0.960537348015+0*(0.02/sqrt(l*w*mult))} lnfactor = 6.14575492391258e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.4667525e-05 lcit = -9.024682925125e-12
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.277998700702905 leta0 = -2.5947385880257e-7
+ etab = -0.02921139354 letab = 2.72689819265577e-8
+ dsub = 0.0588309099500002 ldsub = 4.53057132207125e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.0479946946115999 lpclm = 1.0783082469191e-6
+ pdiblc1 = -0.0068843632690001 lpdiblc1 = 3.79386479565428e-7
+ pdiblc2 = 0.0059964470822665 lpdiblc2 = -4.19168238515769e-9
+ pdiblcb = -0.411701 lpdiblcb = 3.60987317005e-7
+ drout = 1.55012438231795 ldrout = -1.06366824383367e-6
+ pscbe1 = 432633596.7114 lpscbe1 = -124.299268246576
+ pscbe2 = 1.453248063888e-08 lpscbe2 = 2.06195955473267e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -6.3303731508805e-05 lalpha0 = 1.22398274741432e-10 walpha0 = -9.83670105765341e-26 palpha0 = -3.87367706392573e-33
+ alpha1 = 1.933505e-10 lalpha1 = -1.804936585025e-16
+ beta0 = -41.017491252125 lbeta0 = 8.510803942344e-05 pbeta0 = -1.55096364853693e-25
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 6.09038636600001e-09 lagidl = 2.10600000740717e-15
+ bgidl = 782472856.000001 lbgidl = 846.15427105972
+ cgidl = 562.413927750001 lcgidl = -0.000181486373624264
+ egidl = 3.1398290592442 legidl = -2.20386518519396e-6
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.504322175 lkt1 = -1.17320878026625e-7
+ kt2 = -0.019032
+ at = 263567.404 lat = -0.21803633947102
+ ute = -1.343242896 lute = -1.0974014436952e-7
+ ua1 = 5.524e-10
+ ub1 = -3.729725659e-18 lub1 = 1.29594446804797e-25
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.81e-6
+ sbref = 2.81e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.29 pmos
* DC IV MOS Parameters
+ lmin = 8.0e-07 lmax = 1e-06 wmin = 7e-06 wmax = 1.0e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.038439931125+0*(0.0/sqrt(l*w*mult))} lvth0 = 1.9668886054842e-8
+ k1 = 0.5906126265 lk1 = -1.04763779508829e-8
+ k2 = 0.02751640895 lk2 = 7.67582985813028e-9
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 13061.449095 lvsat = 0.0325116929075719
+ ua = -9.06536897720001e-10 lua = 2.4203473270336e-15
+ ub = 3.5868317875e-18 lub = -2.81253087799019e-24
+ uc = 6.3107339585e-12 luc = -6.43763154122954e-18 wuc = -1.23259516440783e-32
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0135845857075 lu0 = 4.04573066162025e-9
+ a0 = 0.712931320600001 la0 = 9.57801142332962e-8
+ keta = -0.15612272205 lketa = 6.66996062872854e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.550106551525001 lags = 1.25439219523654e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0958530090712999+0*(0.009/sqrt(l*w*mult))} lvoff = 1.68938510236889e-8
+ nfactor = {1.77291871495+0*(0.02/sqrt(l*w*mult))} lnfactor = -1.43786575549403e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -1.3337625e-05 lcit = 1.7118264625625e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -1.21860426749999e-05 leta0 = 5.06940288623259e-11
+ etab = 0.00078033929425 letab = -7.28450632878846e-10
+ dsub = 1.5319711835 ldsub = -9.22126678853168e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.04996180999625 lpclm = -7.90538065128049e-7
+ pdiblc1 = 0.18889710180225 lpdiblc1 = 1.9662350301409e-7
+ pdiblc2 = -0.0348197016362825 lpdiblc2 = 3.39103965243514e-08 wpdiblc2 = 2.64697796016969e-23 ppdiblc2 = -2.52435489670724e-29
+ pdiblcb = -0.025
+ drout = 0.333282847401501 ldrout = 7.22594132185118e-8
+ pscbe1 = -69178212.7425003 lpscbe1 = 344.144564937688
+ pscbe2 = 1.840896906885e-08 lpscbe2 = -3.59810173627181e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.00025329086614975 lalpha0 = -1.73144365145817e-10 palpha0 = 7.88860905221012e-31
+ alpha1 = 0.0
+ beta0 = 67.779765317375 lbeta0 = -1.64547435704712e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -2.70605334000001e-09 lagidl = 1.03175204551567e-14
+ bgidl = 1254665040.0 lbgidl = 405.3605063348
+ cgidl = -189.463799999999 lcgidl = 0.000520395244619
+ egidl = 1.87168959037975 legidl = -1.02005065031165e-6
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.580488412500001 lkt1 = -4.6219314489187e-8
+ kt2 = -0.019032
+ at = 48337.625 lat = -0.017118264625625
+ ute = -1.391117025 lute = -6.50494055773772e-8
+ ua1 = 5.524e-10
+ ub1 = -3.5909e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.41e-6
+ sbref = 2.41e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.30 pmos
* DC IV MOS Parameters
+ lmin = 6e-07 lmax = 8.0e-07 wmin = 7e-06 wmax = 1.0e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.946540057525002+0*(0.0/sqrt(l*w*mult))} lvth0 = -4.77401307301255e-8
+ k1 = 0.59524275225 lk1 = -1.38725983391362e-8
+ k2 = 0.0329127025000001 lk2 = 3.71762155773751e-9
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 59860.9299525 lvsat = -0.00181596029880859
+ ua = -2.18776357838e-09 lua = 3.36013350343112e-15
+ ub = 2.580957863135e-18 lub = -2.07471732509884e-24 pub = 1.40129846432482e-45
+ uc = 3.03250253000001e-12 luc = -4.03303239726766e-18
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.00613202721250003 lu0 = 9.51221958049517e-9
+ a0 = 0.94362221325 la0 = -7.34328089799405e-8
+ keta = 0.019410555375 lketa = -6.20549303703394e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = -0.689680622000001 lags = 1.03482931024011e-6
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {0.0153307911677251+0*(0.009/sqrt(l*w*mult))} lvoff = -6.46600223706371e-8
+ nfactor = {1.962272004275+0*(0.02/sqrt(l*w*mult))} lnfactor = -2.82678160035735e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -0.0630409077468501 leta0 = 4.62825765424833e-08 weta0 = 5.45939204284998e-23 peta0 = -8.51969777638693e-29
+ etab = -0.00078033929425 letab = 4.16314915178847e-10
+ dsub = 0.1852475514785 ldsub = 6.57018388527629e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.18595238885375 lpclm = 5.76722165327081e-7
+ pdiblc1 = 0.16298765229625 lpdiblc1 = 2.15628213773989e-7
+ pdiblc2 = 0.02744500370811 lpdiblc2 = -1.17610761692872e-8
+ pdiblcb = -0.025
+ drout = -0.7940560006085 ldrout = 8.99168094928088e-7
+ pscbe1 = 433759236.091001 lpscbe1 = -24.7625684689287
+ pscbe2 = 1.0404743204925e-08 lpscbe2 = 2.2730379560465e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -0.000128252924521375 lalpha0 = 1.06719913030406e-10 walpha0 = -2.06795153138257e-25 palpha0 = -1.97215226305253e-31
+ alpha1 = 0.0
+ beta0 = 25.56667467665 lbeta0 = 1.45087694799539e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 2.42678867225e-08 lagidl = -9.46799945038737e-15
+ bgidl = 2074319252.5 lbgidl = -195.859956805014
+ cgidl = 1293.58225 lcgidl = -0.00056742644828625
+ egidl = -0.281408896629999 legidl = 5.59257855402438e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.7102414755 lkt1 = 4.89552059866273e-8
+ kt2 = -0.019032
+ at = 43672.675 lat = -0.013696500475875
+ ute = -1.6198450625 lute = 1.02723753569065e-7
+ ua1 = 5.53467010000001e-10 lua1 = -7.8265717005015e-19
+ ub1 = -4.3690170425e-18 lub1 = 5.70752741258963e-25
+ uc1 = -2.898021126e-10 luc1 = 1.32472552602663e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.02e-6
+ sbref = 2.01e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.31 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 6e-07 wmin = 7e-06 wmax = 1.0e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.02/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.914622999187028+0*(0.0/sqrt(l*w*mult))} lvth0 = -6.47680409387259e-08 wvth0 = -6.03652813972483e-07 pvth0 = 3.22051794518397e-13
+ k1 = 0.444390559999999 lk1 = 6.66078004872005e-8
+ k2 = 0.0507322538798841 lk2 = -5.78919820118753e-09 wk2 = 1.91935738215305e-08 pk2 = -1.02398676016559e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -2704.27148198453 lvsat = 0.0315628874924961 wvsat = 0.281290277482904 pvsat = -1.50069769488516e-7
+ ua = 1.226709600179e-08 lua = -4.3516063568875e-15 wua = 4.14601084258921e-16 pua = -2.21191751457578e-22
+ ub = -1.25224213060774e-17 lub = 5.98301097857181e-24 wub = 2.38943087821327e-23 pub = -1.27477332068117e-29
+ uc = -1.25620477499999e-12 luc = -1.74498560651362e-18
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0411363862035046 lu0 = -9.16278096300077e-09 wu0 = 1.42310902272595e-08 pu0 = -7.59235779169393e-15
+ a0 = 0.139856216999998 la0 = 3.55380368849416e-7
+ keta = -0.14474227675 lketa = 2.55214263325087e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 1.25
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1246427114985+0*(0.009/sqrt(l*w*mult))} lvoff = 1.00165411693073e-8
+ nfactor = {1.0891138592679+0*(0.02/sqrt(l*w*mult))} lnfactor = 1.8315607611628e-07 wnfactor = -3.04809864056955e-06 pnfactor = 1.62617586523707e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 3.167525e-05 lcit = -1.156385425125e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.00920842325221072 leta0 = 7.73719720782931e-09 weta0 = -1.59227103863488e-06 peta0 = 8.49484560466904e-13
+ etab = 0.0664169194381495 letab = -3.54337586048499e-08 wetab = -3.44619126237054e-07 petab = 1.83856026943099e-13
+ dsub = 0.432939904543 ldsub = -6.6443269968913e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.49935305524623 lpclm = -6.57488657196642e-07 wpclm = -1.06342443276753e-05 ppclm = 5.67342252003642e-12
+ pdiblc1 = 1.751193186706 lpdiblc1 = -6.31687379861285e-7
+ pdiblc2 = 0.00799763922495 lpdiblc2 = -1.38580998069895e-9
+ pdiblcb = -0.025
+ drout = 0.855521778757 ldrout = 1.9110101747696e-8
+ pscbe1 = 494439169.22 lpscbe1 = -57.1356161929161
+ pscbe2 = 1.54395059094e-08 lpscbe2 = -4.13033120604449e-16
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -3.81232336812002e-05 lalpha0 = 5.86352723187186e-11
+ alpha1 = 0.0
+ beta0 = 44.42709312265 lbeta0 = 4.44664193692063e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 2.931681043227e-08 lagidl = -1.21616254941682e-14 wagidl = -2.68511136363387e-13 pagidl = 1.43252033805549e-19
+ bgidl = 2357457500.0 lbgidl = -346.915627537499
+ cgidl = -825.589204953846 lcgidl = 0.000563162118788902 wcgidl = 0.00899810652524417 pcgidl = -4.80053482175039e-9
+ egidl = 1.20727463867 legidl = -2.34962254097788e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.68350575 lkt1 = 3.46915627537504e-8
+ kt2 = -0.019032
+ at = 18000.0
+ ute = -1.665294245 lute = 1.26971119678725e-7
+ ua1 = 5.52e-10
+ ub1 = -8.23768896e-18 lub1 = 2.6347085526048e-24
+ uc1 = -4.1496e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 1.81e-6
+ sbref = 1.81e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.32 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.063267419366+0*(0.0/sqrt(l*w*mult))} wvth0 = 1.42180185466641e-7
+ k1 = 0.59521
+ k2 = 0.02866192842 wk2 = -2.39188007273848e-9
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200000.0
+ ua = 2.7106063484812e-09 wua = -1.36747200730036e-17
+ ub = -3.1082356182e-19 wub = -7.18589113281301e-25
+ uc = -3.9972e-11
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0214334614405 wu0 = -7.06458864340986e-9
+ a0 = 0.911125612687 wa0 = -1.07463754696568e-8
+ keta = -0.0079259
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.119575427913 wags = 7.32940393717753e-9
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.093204657+0*(0.009/sqrt(l*w*mult))}
+ nfactor = {1.65130365316+0*(0.02/sqrt(l*w*mult))} wnfactor = 5.17329490018015e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.08353125
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0029407877
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 333712830.0
+ pscbe2 = 1.5000958e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 5.0667189e-5
+ alpha1 = 0.0
+ beta0 = 38.266046
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -1.23566635609e-08 wagidl = 1.36683986756643e-13
+ bgidl = 1704700000.0
+ cgidl = -39.5608999999999 wcgidl = 0.0051254572987254
+ egidl = 0.69350825
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.57506439519 wkt1 = -4.61291156885278e-9
+ kt2 = -0.019032
+ at = 383654.1836 wat = 0.321195324053459
+ ute = -1.0173591109 wute = -2.55760319206397e-6
+ ua1 = 2.393902706192e-09 wua1 = -1.16939700150493e-14
+ ub1 = -1.8687644069e-18 wub1 = -8.8448308118338e-24
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.33 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.063267419366+0*(0.0/sqrt(l*w*mult))} wvth0 = 1.42180185466641e-7
+ k1 = 0.59521
+ k2 = 0.02866192842 wk2 = -2.39188007273869e-9
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200000.0
+ ua = 2.7106063484812e-09 wua = -1.36747200730036e-17
+ ub = -3.1082356182e-19 wub = -7.18589113281301e-25
+ uc = -3.9972e-11
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0214334614405 wu0 = -7.06458864340991e-9
+ a0 = 0.911125612687 wa0 = -1.07463754696568e-8
+ keta = -0.0079259
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.119575427913 wags = 7.32940393717711e-9
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.093204657+0*(0.009/sqrt(l*w*mult))}
+ nfactor = {1.65130365316+0*(0.02/sqrt(l*w*mult))} wnfactor = 5.17329490018015e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.08353125
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0029407877
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 333712830.0
+ pscbe2 = 1.5000958e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 5.0667189e-5
+ alpha1 = 0.0
+ beta0 = 38.266046
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -1.23566635609e-08 wagidl = 1.36683986756643e-13
+ bgidl = 1704700000.0
+ cgidl = -39.5608999999999 wcgidl = 0.0051254572987254
+ egidl = 0.69350825
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.57506439519 wkt1 = -4.61291156885447e-9
+ kt2 = -0.019032
+ at = 383654.1836 wat = 0.321195324053457
+ ute = -1.0173591109 wute = -2.55760319206397e-6
+ ua1 = 2.393902706192e-09 wua1 = -1.16939700150493e-14
+ ub1 = -1.8687644069e-18 wub1 = -8.84483081183379e-24
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.34 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.06800842414245+0*(0.0/sqrt(l*w*mult))} lvth0 = 3.76127850990202e-08 wvth0 = 1.44280290874126e-07 pvth0 = -1.66611967507977e-14
+ k1 = 0.6042078926875 lk1 = -7.13848266257486e-8
+ k2 = 0.0258520720107467 lk2 = 2.22920098720932e-08 wk2 = 5.37850993494317e-09 pk2 = -6.16464279778928e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 358690.921070056 lvsat = -1.25897521576389 wvsat = -0.418340997170324 pvsat = 3.31891039275575e-6
+ ua = 2.45677234556693e-09 lua = 2.01379333129043e-15 wua = -1.41858017249693e-17 pua = 4.05466884133254e-24
+ ub = 1.20276523993404e-20 lub = -2.5613417222652e-24 wub = -1.14398646462076e-24 pub = 3.37489201383839e-30
+ uc = -5.164762621625e-11 luc = 9.26286389647504e-17
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0207922897795951 lu0 = 5.08673857764685e-09 wu0 = -8.18016463586416e-09 pu0 = 8.85042771401528e-15
+ a0 = 0.94119696678194 la0 = -2.38571238068969e-07 wa0 = -5.24124667540895e-08 pa0 = 3.30558143535494e-13
+ keta = -0.004938304614875 lketa = -2.37021029258661e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.0871268867621089 lags = 2.574306634633e-07 wags = 8.06818856096936e-08 pags = -5.81942280111308e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0947862308566375+0*(0.009/sqrt(l*w*mult))} lvoff = 1.2547424099503e-8
+ nfactor = {1.61132612476985+0*(0.02/sqrt(l*w*mult))} lnfactor = 3.17161921370867e-07 wnfactor = 9.84056915776707e-07 pnfactor = -3.70278436589373e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.652860044042275 lpclm = 5.84216401324086e-06 wpclm = -8.470329472543e-22 ppclm = 3.23117426778526e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00456413311797212 lpdiblc2 = -1.28788189902089e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 563540476.342287 lpscbe1 = -1823.33878139477
+ pscbe2 = -1.55054993344525e-08 lpscbe2 = 2.42023131795166e-13 ppscbe2 = -3.85185988877447e-34
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 7.83237609926249e-05 lalpha0 = -2.1941355218635e-10 walpha0 = -2.06795153138257e-25 palpha0 = -7.88860905221012e-31
+ alpha1 = 0.0
+ beta0 = 39.1457124405462 lbeta0 = -6.9788381044059e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -3.33487714590578e-08 lagidl = 1.66540992970575e-13 wagidl = 2.76401479389901e-13 pagidl = -1.10844942639342e-18
+ bgidl = 1296345515.41866 lbgidl = 3239.6823451985 wbgidl = 1251.662822859 pbgidl = -0.00993007326346601
+ cgidl = -52.7880048261322 lcgidl = 0.000104937302273646 wcgidl = 0.00683914331123034 pcgidl = -1.3595536548638e-8
+ egidl = 1.21251915959209 legidl = -4.11757564630338e-6
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.608220326956748 lkt1 = 2.63042750451153e-07 wkt1 = 1.58859293349513e-07 pkt1 = -1.29690755508087e-12
+ kt2 = -0.019032
+ at = 714488.087097667 lat = -2.62467242756826 wat = -0.276746687564689 pat = 4.74377593888262e-6
+ ute = -0.487574115655178 lute = -4.20305190869978e-06 wute = -5.07268942806387e-06 pute = 1.99534492287364e-11
+ ua1 = 4.72628109065194e-09 lua1 = -1.85039355750049e-14 wua1 = -2.31935423960609e-14 pua1 = 9.12319149826174e-20
+ ub1 = -5.23349222759464e-19 lub1 = -1.06738580904549e-23 wub1 = -1.44411917016906e-23 pub1 = 4.43987571014836e-29
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.35 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.05129232297186+0*(0.0/sqrt(l*w*mult))} lvth0 = -2.81400824360061e-08 wvth0 = 1.93195733521591e-07 pvth0 = -2.09070334981806e-13
+ k1 = 0.6028041533 lk1 = -6.58632107263162e-8
+ k2 = 0.0308769845810631 lk2 = 2.52649115219047e-09 wk2 = -1.27331623638283e-08 pk2 = 9.59592556768576e-15
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -12545.2385325367 lvsat = 0.201284074213703 wvsat = 0.67151370576778 pvsat = -9.68038530524798e-7
+ ua = 3.13468523673447e-09 lua = -6.52780415681577e-16 wua = 9.33765700792385e-16 pua = -3.72471730606823e-21
+ ub = -1.44898058495651e-18 lub = 3.18554148441522e-24 wub = -1.75484210754739e-24 pub = 5.77769573956849e-30
+ uc = -5.52637784975e-11 luc = 1.06852792043809e-16
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0212099025630851 lu0 = 3.44405660572547e-09 wu0 = -5.11422274907537e-09 pu0 = -3.20947002737774e-15
+ a0 = 0.743826641146377 la0 = 5.37785924670145e-07 wa0 = 5.07511899617937e-07 pa0 = -1.8719071512107e-12
+ keta = -0.00501267161000001 lketa = -2.34095799787069e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.0979642604110406 lags = 2.14801800028359e-07 wags = -1.5629825926175e-08 pags = -2.03099681226416e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0637375436500176+0*(0.009/sqrt(l*w*mult))} lvoff = -1.09582742271173e-7
+ nfactor = {1.90494159164811+0*(0.02/sqrt(l*w*mult))} lnfactor = -8.37775985672094e-07 wnfactor = 1.37880798090854e-06 pnfactor = -5.25553965434512e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.0183211905 leta0 = 2.42613905562297e-7
+ etab = -0.12306697823 letab = 2.08739224202596e-7
+ dsub = 0.817977904625 ldsub = -1.01475737773196e-6
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.05151476838812 lpclm = -8.62002833328183e-7
+ pdiblc1 = 0.5839957106185 lpdiblc1 = -7.63083097696422e-7
+ pdiblc2 = -0.00116412829032 lpdiblc2 = 9.65332590061517e-09 ppdiblc2 = 1.26217744835362e-29
+ pdiblcb = 0.1683505 lpdiblcb = -7.605451585025e-07 wpdiblcb = -2.11758236813575e-22 ppdiblcb = 6.05845175209737e-28
+ drout = 0.1346289 ldrout = 1.6731993487055e-6
+ pscbe1 = -159424727.08145 lpscbe1 = 1020.44846109852 ppscbe1 = 8.67361737988404e-19
+ pscbe2 = 7.64564645311875e-08 lpscbe2 = -1.19709712880149e-13
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 4.43365799732225e-05 lalpha0 = -8.57248057106256e-11
+ alpha1 = -9.667525e-11 lalpha1 = 3.8027257925125e-16
+ beta0 = 70.6002512545225 lbeta0 = -0.000130705423801875
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.67527847556901e-08 lagidl = -3.05337289079173e-14 wagidl = -5.22767650783143e-14 pagidl = 1.84408091613529e-19
+ bgidl = 2989897230.66268 lbgidl = -3421.91179447245 wbgidl = -2503.325645718 pbgidl = 0.00484019265262399
+ cgidl = -504.324173199985 lcgidl = 0.00188105707825304 wcgidl = 0.00665313393090154 pcgidl = -1.28638677210678e-8
+ egidl = -1.60756773472605 legidl = 6.97525025293149e-06 wegidl = -1.6940658945086e-21 pegidl = 4.8467614016779e-27
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.5423147225 lkt1 = 3.8027257925123e-09 wkt1 = -1.70848576624177e-7
+ kt2 = -0.019032
+ at = -162530.35277442 lat = 0.825083990760795 wat = 2.58736985724193 pat = -6.52224081069694e-6
+ ute = -1.82569547518022 lute = 1.06045514959879e-06 wute = 8.22538077092878e-07 pute = -3.23545763893523e-12
+ ua1 = -4.9057671776e-10 lua1 = 2.01660069867255e-15 wua1 = -1.97215226305253e-31 pua1 = 2.63310734584192e-36
+ ub1 = -2.65418634019078e-18 lub1 = -2.2921996348532e-24 wub1 = -7.38877964349068e-24 pub1 = 1.66580590084938e-29
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.36 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.16479481403929+0*(0.0/sqrt(l*w*mult))} lvth0 = 1.91317551555322e-07 wvth0 = 5.36607933377802e-07 pvth0 = -8.73059540464782e-13
+ k1 = 0.55879817175 lk1 = 1.92225746305162e-8
+ k2 = 0.0180027216084482 lk2 = 2.74189429810564e-08 wk2 = 6.02546287175858e-08 pk2 = -1.31526333427184e-13
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 132323.17183985 lvsat = -0.0788197215833593 wvsat = 0.330336577145735 pvsat = -3.0837084644843e-7
+ ua = 3.96530972775167e-09 lua = -2.25879702218578e-15 wua = -2.8289005169323e-15 pua = 3.55041663923352e-21
+ ub = 1.63095985574332e-18 lub = -2.7695387573801e-24 wub = -9.97099513799034e-24 pub = 2.16636687046951e-29
+ uc = 5.465298373e-13 luc = -1.05671817306874e-18
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0319904483313898 lu0 = -1.74001825400206e-08 wu0 = -4.26487389484654e-08 pu0 = 6.9363704716724e-14
+ a0 = 1.24657372181402 la0 = -4.34278069536147e-07 wa0 = -1.11171262206291e-06 pa0 = 1.25887155758182e-12
+ keta = 0.04594012976 lketa = -1.21927076191609e-07 pketa = -2.01948391736579e-28
+ a1 = 0.0
+ a2 = 0.5
+ ags = -0.177476008672286 lags = 7.47366937502318e-07 wags = -6.30253763501852e-07 pags = 9.85278775195843e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.256869510875803+0*(0.009/sqrt(l*w*mult))} lvoff = 2.63838882019719e-07 wvoff = 6.69722011790114e-07 pvoff = -1.29491085840625e-12
+ nfactor = {0.424799645578558+0*(0.02/sqrt(l*w*mult))} lnfactor = 2.02408586776312e-06 wnfactor = 3.71287978739174e-06 pnfactor = -9.76847916253942e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.4667525e-05 lcit = -9.024682925125e-12
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.279113373671569 leta0 = -2.61629084560846e-07 weta0 = -7.72513623006226e-09 peta0 = 1.49365895265073e-14
+ etab = -0.02921139354 letab = 2.72689819265577e-8
+ dsub = -0.505373742531682 ldsub = 1.54394964880372e-06 wdsub = 3.91016730878697e-06 pdsub = -7.56032804237615e-12
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.0479946946115986 lpclm = 1.0783082469191e-6
+ pdiblc1 = -0.0068843632690001 lpdiblc1 = 3.79386479565428e-7
+ pdiblc2 = 0.0059964470822665 lpdiblc2 = -4.19168238515769e-9
+ pdiblcb = -0.411701 lpdiblcb = 3.60987317005e-7
+ drout = 1.55012438231795 ldrout = -1.06366824383367e-6
+ pscbe1 = 432633596.7114 lpscbe1 = -124.299268246576
+ pscbe2 = 1.453248063888e-08 lpscbe2 = 2.06195955473267e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -6.3303731508805e-05 lalpha0 = 1.22398274741432e-10 walpha0 = 3.31755453690697e-27 palpha0 = -5.33354700809895e-32
+ alpha1 = 1.933505e-10 lalpha1 = -1.804936585025e-16
+ beta0 = -41.017491252125 lbeta0 = 8.510803942344e-05 pbeta0 = -7.75481824268463e-26
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -3.79933550345672e-09 lagidl = 9.20389837374436e-15 wagidl = 6.85397877824141e-14 pagidl = -4.91913174254535e-20
+ bgidl = 494582812.252974 lbgidl = 1402.79111009481 wbgidl = 1995.19488652466 pbgidl = -0.00385771928906985
+ cgidl = 562.41392775 lcgidl = -0.000181486373624264
+ egidl = 3.1398290592442 legidl = -2.20386518519396e-6
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.45665735173485 lkt1 = -1.61816228868759e-07 wkt1 = -3.30336577145737e-07 pkt1 = 3.0837084644843e-13
+ kt2 = -0.019032
+ at = 482825.59101969 lat = -0.422714953344836 wat = -1.51954825487038 pat = 1.41850589366278e-6
+ ute = -1.10587207613955 lute = -3.31326991563349e-07 wute = -1.64507615418576e-06 pute = 1.53568681531318e-12
+ ua1 = 5.524e-10
+ ub1 = -4.07195909004377e-18 lub1 = 4.49071065851315e-25 wub1 = 2.37181662390637e-24 pub1 = -2.21410267749971e-30
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.81e-6
+ sbref = 2.81e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.37 pmos
* DC IV MOS Parameters
+ lmin = 8.0e-07 lmax = 1e-06 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.702531956385387+0*(0.0/sqrt(l*w*mult))} lvth0 = -2.40207137378885e-07 wvth0 = -2.32797864358327e-06 pvth0 = 1.80104635206124e-12
+ k1 = 0.590612626499999 lk1 = -1.04763779508821e-8
+ k2 = 0.0817000243448977 lk2 = -3.20428076099331e-08 wk2 = -3.75514453234492e-07 pk2 = 2.75266283420491e-13
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 13243.1770870148 lvsat = 0.0323420489183862 wvsat = -0.00125944876622697 pvsat = 1.17570172051707e-9
+ ua = -1.50979324618813e-09 lua = 2.85223897950189e-15 wua = 4.18081141696161e-15 pua = -2.9931844996161e-21
+ ub = -5.71714501715879e-18 lub = 4.08995388199839e-24 wub = 6.44803366708681e-23 pub = -4.78370217955334e-29
+ uc = 6.3107339585e-12 luc = -6.43763154122954e-18 puc = -5.87747175411144e-39
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = -0.0127367446746734 lu0 = 2.43528757671044e-08 wu0 = 1.82417506008596e-07 pu0 = -1.40736760281918e-13
+ a0 = 0.553429650479247 la0 = 2.12775386775221e-07 wa0 = 1.1054113316149e-06 pa0 = -8.10824738796182e-13
+ keta = -0.15612272205 lketa = 6.66996062872853e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.263735352133473 lags = 3.35493926133337e-07 wags = 1.98466867849023e-06 pags = -1.45576439901597e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {0.387323598323788+0*(0.009/sqrt(l*w*mult))} lvoff = -3.37518606383645e-07 wvoff = -3.34861005895056e-06 pvoff = 2.45622222129053e-12
+ nfactor = {6.83062041816155+0*(0.02/sqrt(l*w*mult))} lnfactor = -3.95577985254696e-06 wnfactor = -3.50519262301475e-05 pnfactor = 2.64186610788636e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -1.3337625e-05 lcit = 1.7118264625625e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.000333212278411439 leta0 = -1.38640999952687e-09 weta0 = -2.39375059684739e-09 peta0 = 9.95971438097263e-15
+ etab = -0.0021051576535863 letab = 1.96517519541108e-09 wetab = 1.99976653602664e-08 petab = -1.86679206021355e-14
+ dsub = 4.35302618049806 ldsub = -2.99139097134416e-06 wdsub = -1.95510564775253e-05 pdsub = 1.43408416682653e-11
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.04996180999625 lpclm = -7.90538065128049e-7
+ pdiblc1 = 0.18889710180225 lpdiblc1 = 1.96623503014091e-7
+ pdiblc2 = -0.0348197016362825 lpdiblc2 = 3.39103965243514e-08 wpdiblc2 = 5.29395592033938e-23 ppdiblc2 = -1.26217744835362e-29
+ pdiblcb = -0.025
+ drout = 0.3332828474015 ldrout = 7.22594132185127e-8
+ pscbe1 = -69178212.7424994 lpscbe1 = 344.144564937687
+ pscbe2 = 1.840896906885e-08 lpscbe2 = -3.59810173627181e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.00025329086614975 lalpha0 = -1.73144365145817e-10
+ alpha1 = 0.0
+ beta0 = 67.779765317375 lbeta0 = -1.64547435704711e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 3.49571355826957e-08 lagidl = -2.69754611675345e-14 wagidl = -2.61021190488984e-13 pagidl = 2.58455503595788e-19
+ bgidl = 2694115258.73513 lbgidl = -650.483426358507 wbgidl = -9975.97443262325 pbgidl = 0.00731742712620131
+ cgidl = -189.4638 lcgidl = 0.000520395244619
+ egidl = 1.87168959037975 legidl = -1.02005065031165e-6
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.553364831602275 lkt1 = -7.15393128751184e-08 wkt1 = -1.87977427795077e-07 pkt1 = 1.75477868733843e-13
+ kt2 = -0.019032
+ at = 48337.6250000001 lat = -0.017118264625625
+ ute = -1.391117025 lute = -6.50494055773705e-8
+ ua1 = 5.524e-10
+ ub1 = -3.5909e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.41e-6
+ sbref = 2.41e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.38 pmos
* DC IV MOS Parameters
+ lmin = 6e-07 lmax = 8.0e-07 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.01396927963674+0*(0.0/sqrt(l*w*mult))} lvth0 = -1.17663035873994e-08 wvth0 = 4.67311885498568e-07 pvth0 = -2.49313227472914e-13
+ k1 = 0.59524275225 lk1 = -1.38725983391366e-8
+ k2 = 0.0330392792108561 lk2 = 3.65009224961227e-09 wk2 = -8.77227996377076e-10 pk2 = 4.68005522207034e-16
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 59679.2019604852 lvsat = -0.00171900750642867 wvsat = 0.00125944876622741 pvsat = -6.71922214026011e-10
+ ua = -2.24076305545416e-09 lua = 3.38840898944757e-15 wua = 3.67307893911595e-16 pua = -1.95960597941306e-22
+ ub = 2.97081413257164e-18 lub = -2.28270759412463e-24 wub = -2.70186222884127e-24 pub = 1.44145700839796e-30
+ uc = 3.03250252999999e-12 luc = -4.03303239726765e-18
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0111336155300405 lu0 = 6.84384720514575e-09 wu0 = -3.46630376854124e-08 pu0 = 1.8492903920356e-14
+ a0 = 0.943622213249999 la0 = -7.34328089799413e-8
+ keta = 0.0194105553750001 lketa = -6.20549303703393e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = -0.689680621999999 lags = 1.03482931024011e-6
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {0.0153307911677251+0*(0.009/sqrt(l*w*mult))} lvoff = -6.46600223706371e-8
+ nfactor = {1.4515530583581+0*(0.02/sqrt(l*w*mult))} lnfactor = -1.02070487943387e-08 wnfactor = 3.53948964709615e-06 pnfactor = -1.88833542417403e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -0.0689596709112535 leta0 = 4.94402662845083e-08 weta0 = 4.10194317471605e-08 peta0 = -2.18840719342689e-14
+ etab = 0.00210515765358631 letab = -1.12311213397657e-09 wetab = -1.99976653602665e-08 petab = 1.0668854458029e-14
+ dsub = 0.185215816888849 ldsub = 6.57187694150145e-08 wdsub = 2.19933590518131e-10 pdsub = -1.1733567021053e-16
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.18595238885375 lpclm = 5.76722165327082e-7
+ pdiblc1 = 0.16298765229625 lpdiblc1 = 2.15628213773989e-7
+ pdiblc2 = 0.02744500370811 lpdiblc2 = -1.17610761692872e-8
+ pdiblcb = -0.025
+ drout = -0.794056000608499 ldrout = 8.99168094928088e-7
+ pscbe1 = 433759236.091 lpscbe1 = -24.7625684689292
+ pscbe2 = 1.0404743204925e-08 lpscbe2 = 2.27303795604648e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -0.000128252924521375 lalpha0 = 1.06719913030406e-10 palpha0 = 1.97215226305253e-31
+ alpha1 = 0.0
+ beta0 = 25.56667467665 lbeta0 = 1.45087694799539e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -2.4066334437246e-08 lagidl = 1.63185492094429e-14 wagidl = 3.3497577633083e-13 pagidl = -1.7871125155138e-19
+ bgidl = 2074319252.5 lbgidl = -195.859956805012
+ cgidl = 1293.58225 lcgidl = -0.00056742644828625
+ egidl = -0.281408896629999 legidl = 5.59257855402438e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.737365056397725 lkt1 = 6.34257720134687e-08 wkt1 = 1.87977427795077e-07 pkt1 = -1.00286897615813e-13
+ kt2 = -0.019032
+ at = 43672.675 lat = -0.013696500475875
+ ute = -1.6198450625 lute = 1.02723753569061e-7
+ ua1 = 5.5346701e-10 lua1 = -7.8265717005015e-19
+ ub1 = -4.3690170425e-18 lub1 = 5.70752741258963e-25
+ uc1 = -2.898021126e-10 luc1 = 1.32472552602663e-16 wuc1 = -7.88860905221012e-31
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.02e-6
+ sbref = 2.01e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.39 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 6e-07 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.14638131499707+0*(0.0/sqrt(l*w*mult))} lvth0 = 5.88761793375101e-08 wvth0 = 1.00252640846733e-06 pvth0 = -5.3485285154936e-13
+ k1 = 0.319675857645699 lk1 = 1.33143717766731e-07 wk1 = 8.64323521484468e-07 pk1 = -4.61120920329571e-13
+ k2 = 0.0558314447618026 lk2 = -8.50964203264554e-09 wk2 = -1.61458892616629e-08 pk2 = 8.61391265054358e-15
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 104666.324331749 lvsat = -0.0257198622271097 wvsat = -0.462831543968169 pvsat = 2.46922942864738e-7
+ ua = 1.89201604729619e-08 lua = -7.90104951758005e-15 wua = -4.56938368451374e-14 pua = 2.4377890426065e-20
+ ub = -9.96242176075601e-18 lub = 4.61723842114514e-24 wub = 6.15247257324026e-24 pub = -3.28237488018656e-30
+ uc = -5.00541716893279e-11 luc = 2.42889737321149e-17 wuc = 3.3818972269086e-16 puc = -1.80425908004187e-22
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.067808945364426 lu0 = -2.33927246381481e-08 wu0 = -1.70620573816945e-07 pu0 = 9.10269292342091e-14
+ a0 = -1.57868459581877 la0 = 1.27223048519229e-06 wa0 = 1.19101855604041e-05 pa0 = -6.35414354740339e-12
+ keta = -0.0354592822105759 lketa = -3.27815976692465e-08 wketa = -7.57375521053992e-07 pketa = 4.0406362735991e-13
+ a1 = 0.0
+ a2 = 0.5
+ ags = 1.25
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.460411666489074+0*(0.009/sqrt(l*w*mult))} lvoff = 1.89150957501554e-07 wvoff = 2.32701518028041e-06 pvoff = -1.2414742337555e-12
+ nfactor = {-2.44847786316903+0*(0.02/sqrt(l*w*mult))} lnfactor = 2.070478947995e-06 wnfactor = 2.14688482581577e-05 pnfactor = -1.14537378899684e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 3.167525e-05 lcit = -1.156385425125e-11 wcit = -1.03397576569128e-25
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -0.645107384117879 leta0 = 3.56817952018809e-07 weta0 = 2.94240315865763e-06 peta0 = -1.56978679715964e-12
+ etab = -0.0514765095049123 letab = 2.74629752034183e-08 wetab = 4.72430201070515e-07 petab = -2.52043874422125e-13
+ dsub = 0.548560692932572 ldsub = -1.28127538678692e-07 wdsub = -8.01299005579815e-07 pdsub = 4.2749702597186e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.664173587097295 lpclm = 1.03026862412684e-06 wpclm = 1.12902796955821e-05 ppclm = -6.02342066899153e-12
+ pdiblc1 = 2.80557039401771 lpdiblc1 = -1.19420289184812e-06 wpdiblc1 = -7.3072621238163e-06 ppdiblc1 = 3.89846087936662e-12
+ pdiblc2 = 0.0418571444378737 lpdiblc2 = -1.94500253093198e-08 wpdiblc2 = -2.34660118084678e-07 ppdiblc2 = 1.25192346298766e-13
+ pdiblcb = -0.025
+ drout = -1.03539131722172 ldrout = 1.02792169301783e-06 wdrout = 1.31047954658496e-05 pdrout = -6.99147390500806e-12
+ pscbe1 = 12924466.5882235 lpscbe1 = 199.75488523465 wpscbe1 = 3337.09238420748 ppscbe1 = -0.00178035547243661
+ pscbe2 = 1.51456515674432e-08 lpscbe2 = -2.562603598988e-16 wpscbe2 = 2.03652989462365e-15 ppscbe2 = -1.08649888143114e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -0.000605098766252098 lalpha0 = 3.61119553822956e-10 walpha0 = 3.92937063278255e-09 palpha0 = -2.09633887944265e-15
+ alpha1 = 0.0
+ beta0 = 0.0719191629364104 lbeta0 = 2.81103490202977e-05 wbeta0 = 0.000307399363741443 pbeta0 = -1.63999097552879e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 5.89772458722511e-09 lagidl = 3.32573899592472e-16 wagidl = -1.06207363308373e-13 pagidl = 5.66621593618336e-20
+ bgidl = 3582162289.18619 lbgidl = -1000.30175609228 wbgidl = -8487.70141920471 pbgidl = 0.00452823114565282
+ cgidl = 2887.9746879239 lcgidl = -0.00141804278588084 wcgidl = -0.0167383989593391 pcgidl = 8.93001953680222e-9
+ egidl = 1.30409385745434 legidl = -2.8661579141533e-07 wegidl = -6.70996494778341e-07 pegidl = 3.57979984946712e-13
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.469770184696999 lkt1 = -7.93374300132271e-08 wkt1 = -1.4812742441893e-06 pkt1 = 7.90267215646215e-13
+ kt2 = -0.019032
+ at = 18000.0
+ ute = -1.665294245 lute = 1.26971119678726e-7
+ ua1 = 5.52e-10
+ ub1 = -1.60817842066201e-17 lub1 = 6.81957258715286e-24 wub1 = 5.43627647617475e-23 pub1 = -2.90028068142161e-29
+ uc1 = -4.1496e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 1.81e-6
+ sbref = 1.81e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.40 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.054497420288+0*(0.0/sqrt(l*w*mult))} wvth0 = 9.89405293924761e-8
+ k1 = 0.59521
+ k2 = 0.0295483765283 wk2 = -6.76242914458949e-9
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200000.0
+ ua = 2.7074193197134e-09 wua = 2.03862568593801e-18
+ ub = -3.4487757531e-19 wub = -5.50689000846123e-25
+ uc = -3.9972e-11
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0211469748272 wu0 = -5.65209332627584e-9
+ a0 = 0.909778235304 wa0 = -4.10325793625426e-9
+ keta = -0.0079259
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.1122159834078 wags = 4.36144532822825e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.093204657+0*(0.009/sqrt(l*w*mult))}
+ nfactor = {1.78357068798+0*(0.02/sqrt(l*w*mult))} wnfactor = -1.34800692060718e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.08353125
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0029407877
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 333712830.0
+ pscbe2 = 1.5000958e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 5.0667189e-5
+ alpha1 = 0.0
+ beta0 = 38.266046
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.6231934973e-08 wagidl = -4.26941098648905e-15
+ bgidl = 1600670587 wbgidl = 512.907242031677
+ cgidl = 1000.0
+ egidl = 0.69350825
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.576
+ kt2 = -0.019032
+ at = 448800.0
+ ute = -1.5361
+ ua1 = 2.2096e-11
+ ub1 = -3.6627e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.41 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.054497420288+0*(0.0/sqrt(l*w*mult))} wvth0 = 9.89405293924761e-8
+ k1 = 0.59521
+ k2 = 0.0295483765283 wk2 = -6.76242914458944e-9
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200000.0
+ ua = 2.7074193197134e-09 wua = 2.03862568593485e-18
+ ub = -3.4487757531e-19 wub = -5.50689000846123e-25
+ uc = -3.9972e-11
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0211469748272 wu0 = -5.65209332627584e-9
+ a0 = 0.909778235304 wa0 = -4.10325793625257e-9
+ keta = -0.0079259
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.1122159834078 wags = 4.36144532822823e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.093204657+0*(0.009/sqrt(l*w*mult))}
+ nfactor = {1.78357068798+0*(0.02/sqrt(l*w*mult))} wnfactor = -1.34800692060718e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.08353125
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0029407877
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 333712830.0
+ pscbe2 = 1.5000958e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 5.0667189e-5
+ alpha1 = 0.0
+ beta0 = 38.266046
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.6231934973e-08 wagidl = -4.26941098648902e-15
+ bgidl = 1600670587 wbgidl = 512.907242031677
+ cgidl = 1000.0
+ egidl = 0.69350825
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.576
+ kt2 = -0.019032
+ at = 448800.0
+ ute = -1.5361
+ ua1 = 2.2096e-11
+ ub1 = -3.6627e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.42 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.05693937569188+0*(0.0/sqrt(l*w*mult))} lvth0 = 1.93732654064793e-08 wvth0 = 8.97053879791374e-08 pvth0 = 7.3267040578442e-14
+ k1 = 0.6042078926875 lk1 = -7.13848266257453e-8
+ k2 = 0.0283445039407229 lk2 = 9.5509291929061e-09 wk2 = -6.91019140720289e-09 pk2 = 1.17227264925487e-15
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 273841.7226125 lvsat = -0.585823675554882
+ ua = 2.44989507539687e-09 lua = 2.04306987990643e-15 wua = 1.97219323850995e-17 pua = -1.40290602114341e-22
+ ub = -1.9497362761997e-19 lub = -1.18926371851859e-24 wub = -1.23386111605879e-25 pub = -3.39000960830193e-30
+ uc = -5.164762621625e-11 luc = 9.26286389647506e-17
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0200674461306593 lu0 = 8.56444631164957e-09 wu0 = -4.60639116008856e-09 pu0 = -8.29608336395743e-15
+ a0 = 0.927987831199286 la0 = -1.44465920083223e-07 wa0 = 1.27139345774357e-08 pa0 = -1.3341928089332e-13
+ keta = -0.004938304614875 lketa = -2.37021029258661e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.0891245598534977 lags = 1.83195924225175e-07 wags = 7.08325462138711e-08 pags = -2.15934876363223e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0947862308566376+0*(0.009/sqrt(l*w*mult))} lvoff = 1.2547424099503e-8
+ nfactor = {1.89891585075407+0*(0.02/sqrt(l*w*mult))} lnfactor = -9.15091425593903e-07 wnfactor = -4.3387719475422e-07 pnfactor = 2.37272492950142e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.652860044042275 lpclm = 5.84216401324086e-06 wpclm = 4.2351647362715e-22 ppclm = -1.61558713389263e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00456413311797213 lpdiblc2 = -1.28788189902089e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 563540476.342288 lpscbe1 = -1823.33878139477
+ pscbe2 = -1.55054993344525e-08 lpscbe2 = 2.42023131795166e-13 ppscbe2 = 9.62964972193618e-35
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 7.8323760992625e-05 lalpha0 = -2.1941355218635e-10
+ alpha1 = 0.0
+ beta0 = 39.1457124405463 lbeta0 = -6.9788381044059e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 2.65963275777622e-08 lagidl = -8.22259605518442e-14 wagidl = -1.91521965718308e-14 pagidl = 1.18072653855237e-19
+ bgidl = 1343882124.07936 lbgidl = 2037.23255452322 wbgidl = 1017.28804229863 pbgidl = -0.00400150760082188
+ cgidl = 1334.347925 lcgidl = -0.00265255093472713
+ egidl = 1.21251915959209 legidl = -4.11757564630338e-06 pegidl = 6.46234853557053e-27
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.576
+ kt2 = -0.019032
+ at = 649654.770051962 lat = -1.59348232248109 wat = 0.0429078877973579 pat = -3.40409942379776e-7
+ ute = -1.516432475 lute = -1.56032407925125e-7
+ ua1 = 2.2096e-11
+ ub1 = -3.27513178283466e-18 lub1 = -3.07477438872228e-24 wub1 = -8.73786456800493e-25 pub1 = 6.93218922395903e-30
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.43 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.03078803890709+0*(0.0/sqrt(l*w*mult))} lvth0 = -8.34931485931868e-08 wvth0 = 9.21012883429289e-08 pvth0 = 6.38427545179614e-14
+ k1 = 0.6028041533 lk1 = -6.58632107263162e-8
+ k2 = 0.0287548750134528 lk2 = 7.93673252646751e-09 wk2 = -2.27030061902471e-09 pk2 = -1.70787609654978e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 137818.108382575 lvsat = -0.0507741088634006 wvsat = -0.0698386420425674 pvsat = 2.7471064766765e-7
+ ua = 3.40502193217877e-09 lua = -1.71392638687948e-15 wua = -3.9910396444638e-16 pua = 1.50716315720176e-21
+ ub = -1.6318644351322e-18 lub = 4.4627534572848e-24 wub = -8.53150475338072e-25 pub = -5.19477834739526e-31
+ uc = -5.52637784975e-11 luc = 1.06852792043809e-16
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0219128754706398 lu0 = 1.30544077568954e-09 wu0 = -8.58016459032029e-09 pu0 = 7.3347742927262e-15
+ a0 = 0.892998561458087 la0 = -6.83545260987044e-09 wa0 = -2.27966231318439e-07 pa0 = 8.13297355058937e-13
+ keta = -0.00501267161000001 lketa = -2.34095799787069e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.0968820241888725 lags = 1.52681899474657e-07 wags = -1.02939619629796e-08 pags = 1.03176649182958e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0637375436500175+0*(0.009/sqrt(l*w*mult))} lvoff = -1.09582742271173e-7
+ nfactor = {2.13287662828649+0*(0.02/sqrt(l*w*mult))} lnfactor = -1.83537731382154e-06 wnfactor = 2.54995708656491e-07 pnfactor = -3.36960080429135e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.0183211905 leta0 = 2.42613905562297e-7
+ etab = -0.12306697823 letab = 2.08739224202596e-7
+ dsub = 0.817977904625 ldsub = -1.01475737773196e-6
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.05151360686742 lpclm = -8.61998264480684e-07 wpclm = 5.72676864832528e-12 ppclm = -2.25262731077813e-17
+ pdiblc1 = 0.5839957106185 lpdiblc1 = -7.63083097696423e-7
+ pdiblc2 = -0.00116412829032 lpdiblc2 = 9.65332590061517e-09 ppdiblc2 = 6.31088724176809e-30
+ pdiblcb = 0.1683505 lpdiblcb = -7.605451585025e-07 wpdiblcb = 5.29395592033938e-23 ppdiblcb = 3.02922587604869e-28
+ drout = 0.1346289 ldrout = 1.6731993487055e-6
+ pscbe1 = -159424727.08145 lpscbe1 = 1020.44846109852
+ pscbe2 = 7.64564645311875e-08 lpscbe2 = -1.19709712880149e-13
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 4.43365799732225e-05 lalpha0 = -8.57248057106256e-11
+ alpha1 = -9.667525e-11 lalpha1 = 3.8027257925125e-16
+ beta0 = 70.6002512545225 lbeta0 = -0.000130705423801876
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.26604812275049e-09 lagidl = 1.74108203358418e-14 wagidl = 2.40791341371509e-14 pagidl = -5.1978001645196e-20
+ bgidl = 2482165079.25 lbgidl = -2440.20914105527 wbgidl = 3.63797880709171e-12
+ cgidl = 845.084766125 lcgidl = -0.000728031852976518
+ egidl = -1.60756773472605 legidl = 6.97525025293149e-06 wegidl = -4.2351647362715e-22 pegidl = 8.07793566946316e-28
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.5769667525 lkt1 = 3.80272579251315e-9
+ kt2 = -0.019032
+ at = 474458.9061279 lat = -0.904348515756474 wat = -0.553245806785621 pat = 2.00456359603084e-6
+ ute = -1.65886579075 lute = 4.04229751744078e-7
+ ua1 = -4.9057671776e-10 lua1 = 2.01660069867255e-15 pua1 = -1.22251412485518e-36
+ ub1 = -5.25926309515408e-18 lub1 = 4.7298160489427e-24 wub1 = 5.45530641964091e-24 pub1 = -1.79633292509876e-29
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.44 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.04152659863678+0*(0.0/sqrt(l*w*mult))} lvth0 = -6.27300896630299e-08 wvth0 = -7.11544154520299e-08 pvth0 = 3.79498474084032e-13
+ k1 = 0.55879817175 lk1 = 1.92225746305158e-8
+ k2 = 0.0389267126181375 lk2 = -1.17305663413783e-08 wk2 = -4.2909142100532e-08 pk2 = 6.14966422332037e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 170993.27183985 lvsat = -0.114918453283859 wvsat = 0.139677284085135 pvsat = -1.30389443079894e-7
+ ua = 3.16029648891213e-09 lua = -1.24074851869621e-15 wua = 1.14014158592159e-15 pua = -1.46897581066244e-21
+ ub = -1.1603484364625e-18 lub = 3.55107491627695e-24 wub = 3.791288013751e-24 pub = -9.49952287558569e-30
+ uc = 5.465298373e-13 luc = -1.05671817306874e-18
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0211996492725841 lu0 = 2.68446719576116e-09 wu0 = 1.05542814758648e-08 pu0 = -2.96617728484728e-14
+ a0 = 0.968591622029884 la0 = -1.52995013190744e-07 wa0 = 2.58851990605392e-07 pa0 = -1.27968111121901e-13
+ keta = 0.04594012976 lketa = -1.21927076191609e-07 pketa = -2.52435489670724e-29
+ a1 = 0.0
+ a2 = 0.5
+ ags = -0.371631075074579 lags = 1.05855431946604e-06 wags = 3.27009540818412e-07 pags = -5.49001359962375e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0635988679177671+0*(0.009/sqrt(l*w*mult))} lvoff = -1.09850872492858e-07 wvoff = -2.83180725874043e-07 pvoff = 5.47531349381092e-13
+ nfactor = {1.69001496723262+0*(0.02/sqrt(l*w*mult))} lnfactor = -9.79102077865587e-07 wnfactor = -2.52514542578339e-06 pnfactor = 5.03845670371604e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.4667525e-05 lcit = -9.024682925125e-12
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.28882850138512 leta0 = -2.80413332570636e-07 weta0 = -5.56246601997219e-08 peta0 = 1.07550558619463e-13
+ etab = -0.02921139354 letab = 2.72689819265577e-8
+ dsub = 0.287697646912837 ldsub = 1.05421519557952e-08 wdsub = 3.3718413735488e-12 pdsub = -6.51947215364239e-18
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.047997017653008 lpclm = 1.07830607834833e-06 wpclm = -1.14535372949565e-11 ppclm = 1.06919343328136e-17
+ pdiblc1 = -0.00688436326899999 lpdiblc1 = 3.79386479565428e-7
+ pdiblc2 = 0.0059964470822665 lpdiblc2 = -4.19168238515769e-9
+ pdiblcb = -0.411701 lpdiblcb = 3.60987317005e-7
+ drout = 1.55012438231795 ldrout = -1.06366824383367e-6
+ pscbe1 = 432633596.7114 lpscbe1 = -124.299268246576
+ pscbe2 = 1.453248063888e-08 lpscbe2 = 2.06195955473267e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -6.3303731508805e-05 lalpha0 = 1.22398274741432e-10 walpha0 = -3.45323861260498e-27 palpha0 = -3.03525806919044e-32
+ alpha1 = 1.933505e-10 lalpha1 = -1.804936585025e-16
+ beta0 = -41.017491252125 lbeta0 = 8.510803942344e-05 pbeta0 = -5.16987882845642e-26
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 6.74346840257747e-09 lagidl = 6.8202008376949e-15 wagidl = 1.65594841472796e-14 pagidl = -3.743872079153e-20
+ bgidl = 899254331.5 lbgidl = 620.356704273093
+ cgidl = 1317.42535598628 lcgidl = -0.00164130474517625 wcgidl = -0.00372251287584473 pcgidl = 7.19749725801016e-9
+ egidl = 3.1398290592442 legidl = -2.20386518519396e-6
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.523657225 lkt1 = -9.92715121763752e-8
+ kt2 = -0.019032
+ at = -14984.998463649 lat = 0.0419937209908086 wat = 0.93486006238181 pat = -8.72696542533731e-7
+ ute = -1.439531445 lute = -1.9854302435275e-8
+ ua1 = 5.524e-10
+ ub1 = -2.08687233735319e-18 lub1 = -1.40401734321911e-24 wub1 = -7.41546701207983e-24 pub1 = 6.92237553311158e-30
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.81e-6
+ sbref = 2.81e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.45 pmos
* DC IV MOS Parameters
+ lmin = 8.0e-07 lmax = 1e-06 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.49219430894229+0*(0.0/sqrt(l*w*mult))} lvth0 = 3.57970471245718e-07 wvth0 = 1.56537735743742e-06 pvth0 = -1.14821211856713e-12
+ k1 = 0.5906126265 lk1 = -1.04763779508829e-8
+ k2 = -0.0162063490689196 lk2 = 3.97364224087978e-08 wk2 = 1.07203717683233e-07 pk2 = -7.863446293924e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 12987.7318424999 lvsat = 0.0325805083313671
+ ua = -2.51468654978967e-10 lua = 1.94415130195185e-15 wua = -2.02323969748359e-15 pua = 1.48405643430269e-21
+ ub = 1.34054220619851e-17 lub = -1.00461446728764e-23 wub = -2.98016827915453e-23 pub = 2.18596833360124e-29
+ uc = 6.3107339585e-12 luc = -6.43763154122954e-18 puc = 2.93873587705572e-39
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0443506427748238 lu0 = -1.89271009935471e-08 wu0 = -9.90464915967288e-08 pu0 = 7.26510968186586e-14
+ a0 = 0.662356531911316 la0 = 1.3287697461039e-07 wa0 = 5.6835758184093e-07 pa0 = -4.16893128068232e-13
+ keta = -0.15612272205 lketa = 6.66996062872853e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.913448635642713 lags = -1.41074015887107e-07 wags = -1.21868159280342e-06 pags = 8.93909041729269e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.57902961646639+0*(0.009/sqrt(l*w*mult))} lvoff = 3.71306308431024e-07 wvoff = 1.41590362937022e-06 pvoff = -1.0385723916612e-12
+ nfactor = {-2.9977852638955+0*(0.02/sqrt(l*w*mult))} lnfactor = 3.39698287689367e-06 wnfactor = 1.34061041151006e-05 pnfactor = -9.83344439894686e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -1.3337625e-05 lcit = 1.7118264625625e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -0.056562112689848 leta0 = 4.2010532621417e-08 weta0 = 2.78123300998609e-07 peta0 = -2.04004831898985e-13
+ etab = 0.001950829898 letab = -1.82110946393249e-9
+ dsub = 0.387624625673066 ldsub = -8.27401823517723e-08 wdsub = -1.68592068643559e-11 pdsub = 1.23663125306434e-17
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.04996180999625 lpclm = -7.90538065128049e-7
+ pdiblc1 = 0.18889710180225 lpdiblc1 = 1.96623503014091e-7
+ pdiblc2 = -0.0348197016362825 lpdiblc2 = 3.39103965243514e-08 wpdiblc2 = 1.98523347012727e-23 ppdiblc2 = 1.89326617253043e-29
+ pdiblcb = -0.025
+ drout = 0.3332828474015 ldrout = 7.22594132185135e-8
+ pscbe1 = -69178212.7425003 lpscbe1 = 344.144564937687
+ pscbe2 = 1.840896906885e-08 lpscbe2 = -3.59810173627184e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.00025329086614975 lalpha0 = -1.73144365145817e-10
+ alpha1 = 0.0
+ beta0 = 67.7797653173751 lbeta0 = -1.64547435704711e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 4.306638894215e-09 lagidl = 9.09499336789886e-15 wagidl = -1.09901797713119e-13 pagidl = 8.06135181315611e-20
+ bgidl = 670757662.5 lbgidl = 833.659487267938
+ cgidl = -3964.5209411814 lcgidl = 0.00328941853296127 wcgidl = 0.0186125643792236 pcgidl = -1.36524090349824e-8
+ egidl = 1.87168959037975 legidl = -1.02005065031165e-6
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.5914909875 lkt1 = -3.59483557138126e-8
+ kt2 = -0.019032
+ at = 48337.6250000001 lat = -0.017118264625625
+ ute = -1.391117025 lute = -6.50494055773738e-8
+ ua1 = 5.524e-10
+ ub1 = -3.5909e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.41e-6
+ sbref = 2.41e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.46 pmos
* DC IV MOS Parameters
+ lmin = 6e-07 lmax = 8.0e-07 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.763708893211167+0*(0.0/sqrt(l*w*mult))} lvth0 = -1.76377223620144e-07 wvth0 = -7.66573425296422e-07 pvth0 = 5.62285440322055e-13
+ k1 = 0.622953773584957 lk1 = -3.41987710434341e-08 wk1 = -1.36626585856e-07 pk1 = 1.00216283858306e-13
+ k2 = 0.0327284693184924 lk2 = 3.84248844753919e-09 wk2 = 6.55190961791859e-10 pk2 = -4.8058584642915e-16
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 126588.838409808 lvsat = -0.0507464713412859 wvsat = -0.32863222424133 pvsat = 2.41053379642137e-7
+ ua = -8.89625620971965e-09 lua = 8.28514619729192e-15 wua = 3.31815912746611e-14 pua = -2.43388631079203e-20
+ ub = 5.58877062254782e-18 lub = -4.31259175879194e-24 wub = -1.56094506147588e-23 pub = 1.14496100731786e-29
+ uc = 1.10886318918636e-11 luc = -9.94224356484141e-18 wuc = -3.97199885425084e-17 puc = 2.91348101958727e-23
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = -0.0215836746013462 lu0 = 2.94360504734604e-08 wu0 = 1.26646485882117e-07 pu0 = -9.28958306269623e-14
+ a0 = 1.09030692844054 la0 = -1.81026780995778e-07 wa0 = -7.23215199883727e-07 pa0 = 5.30481965190714e-13
+ keta = 0.229998683658141 lketa = -2.16522375406665e-07 wketa = -1.03828497121597e-06 pketa = 7.61587217811769e-13
+ a1 = 0.0
+ a2 = 0.5
+ ags = -2.75678992575627 lags = 2.55106432009185e-06 wags = 1.01916881138957e-05 pags = -7.47565418998308e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {0.144491545024242+0*(0.009/sqrt(l*w*mult))} lvoff = -1.59400081128162e-07 wvoff = -6.36814955778696e-07 pvoff = 4.67106954138452e-13
+ nfactor = {2.92357769181471+0*(0.02/sqrt(l*w*mult))} lnfactor = -9.46366457934553e-07 wnfactor = -3.71818943784614e-06 pnfactor = 2.72731054360733e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -0.152368038034247 leta0 = 1.1228465789116e-07 weta0 = 4.52256545460571e-07 peta0 = -3.31732437378056e-13
+ etab = -0.001950829898 letab = 1.04077750473249e-9
+ dsub = 0.0540186042002024 ldsub = 1.6196150242868e-07 wdsub = 6.47075458213903e-07 pdsub = -4.74633083977188e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.966061993649285 lpclm = 1.42173047496497e-06 wpclm = 5.67989862357925e-06 ppclm = -4.1662340398885e-12
+ pdiblc1 = -0.267737572080258 lpdiblc1 = 5.31567319480279e-07 wpdiblc1 = 2.12365023061728e-06 ppdiblc1 = -1.55770806240893e-12
+ pdiblc2 = 0.0509381824682659 lpdiblc2 = -2.89934402557554e-08 wpdiblc2 = -1.15830909518145e-07 ppdiblc2 = 8.49625512861071e-14
+ pdiblcb = -0.025
+ drout = -2.59017707707413 ldrout = 2.21663188512101e-06 wdrout = 8.85560613213258e-06 pdrout = -6.49563137594991e-12
+ pscbe1 = 483223370.089242 lpscbe1 = -61.0447580773091 wpscbe1 = -243.878263049734 ppscbe1 = 0.000178885925338295
+ pscbe2 = 5.86426695416572e-09 lpscbe2 = 5.60349998835968e-15 wpscbe2 = 2.2386391349601e-14 ppscbe2 = -1.64205299868891e-20
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -0.00034142984455858 lalpha0 = 2.63086249762297e-10 walpha0 = 1.05104876561296e-09 palpha0 = -7.70949524820932e-16
+ alpha1 = 0.0
+ beta0 = -3.41512172328839 lbeta0 = 3.57670620482907e-05 wbeta0 = 0.000142892022861035 pbeta0 = -1.04812013228683e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 6.40925772432472e-08 lagidl = -3.47582913408081e-14 wagidl = -9.96834507721434e-14 pagidl = 7.3118309558621e-20
+ bgidl = 2465556662.32076 lbgidl = -482.834553095588 wbgidl = -1928.95927280472 pbgidl = 0.00141490127139863
+ cgidl = 2427.03728344675 lcgidl = -0.00139882138259461 wcgidl = -0.00558839349763606 pcgidl = 4.09911457248354e-9
+ egidl = -1.39854686775388 legidl = 1.37868414291166e-06 wegidl = 5.50794375565699e-06 pegidl = -4.04010428449318e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.804767472579525 lkt1 = 1.20491012474445e-07 wkt1 = 5.20298704952322e-07 pkt1 = -3.81641701576054e-13
+ kt2 = -0.019032
+ at = 43672.675 lat = -0.013696500475875
+ ute = -1.73709903147725 lute = 1.88730126083721e-07 wute = 5.78109672169248e-07 pute = -4.24046335084504e-13
+ ua1 = 5.5346701e-10 lua1 = -7.82657170049756e-19
+ ub1 = -4.3690170425e-18 lub1 = 5.70752741258963e-25
+ uc1 = -2.898021126e-10 luc1 = 1.32472552602663e-16 wuc1 = 3.94430452610506e-31
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.02e-6
+ sbref = 2.01e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.47 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 6e-07 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.02/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.16431697022375+0*(0.0/sqrt(l*w*mult))} lvth0 = 3.73491885064552e-08 wvth0 = 1.09095647061087e-06 pvth0 = -4.28716046793967e-13
+ k1 = 0.327577581515492 lk1 = 1.23385904306586e-07 wk1 = 8.25364814706486e-07 pk1 = -4.13010938298784e-13
+ k2 = 0.0739546618011692 lk2 = -1.81518913729312e-08 wk2 = -1.05500707291858e-07 pk2 = 5.61541166513843e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 318751.665774059 lvsat = -0.153266300554251 wvsat = -1.51835919592738 pvsat = 8.75778667671504e-7
+ ua = 2.20384300678177e-08 lua = -8.21866360520567e-15 wua = -6.1068171965232e-14 pua = 2.59438568293789e-20
+ ub = -1.58206200025521e-17 lub = 7.109425186652e-24 wub = 3.50357683337812e-23 pub = -1.55698674619622e-29
+ uc = -1.63686061297409e-10 luc = 8.33009291251016e-17 wuc = 8.98441073005881e-16 puc = -4.71378806945501e-22
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0728442822100031 lu0 = -2.09417366251784e-08 wu0 = -1.95446828812399e-07 pu0 = 7.89425632291355e-14
+ a0 = 1.34983104581441 la0 = -3.19484195235324e-07 wa0 = -2.52858553019799e-06 pa0 = 1.49365606326503e-12
+ keta = -0.135501782963306 lketa = -2.15260489617895e-08 wketa = -2.64125375087725e-07 pketa = 3.4856920247937e-13
+ a1 = 0.0
+ a2 = 0.5
+ ags = -1.34861335354646 lags = 1.79979507793506e-06 wags = 1.28122188700056e-05 pags = -8.87372045102148e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.167093472266216+0*(0.009/sqrt(l*w*mult))} lvoff = 6.83208352138414e-09 wvoff = 8.80837395574859e-07 pvoff = -3.42568163570426e-13
+ nfactor = {0.0271341156643778+0*(0.02/sqrt(l*w*mult))} lnfactor = 5.98900672159535e-07 wnfactor = 9.26307610404557e-06 pnfactor = -4.1982595293196e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 6.34338913257499e-05 lcit = -2.85072481917442e-11 wcit = -1.56582995744325e-10 pcit = 8.35378111445764e-17
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.792368295026858 leta0 = -3.91736899478605e-07 weta0 = -4.14493555465166e-06 peta0 = 2.12089253399232e-12
+ etab = 0.0133531442443332 letab = -7.12396922007298e-09 wetab = 1.52793687247313e-07 petab = -8.15161961148776e-14
+ dsub = 0.665424053749745 ldsub = -1.64226361933248e-07 wdsub = -1.37748282093297e-06 pdsub = 6.05478880739066e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.255296675985267 lpclm = 7.70129517921589e-07 wpclm = 6.75691799365828e-06 ppclm = -4.74082925892251e-12
+ pdiblc1 = 0.893254833691984 lpdiblc1 = -8.78279339612403e-08 wpdiblc1 = 2.12122998870702e-06 ppdiblc1 = -1.55641685124859e-12
+ pdiblc2 = -0.079024355704854 lpdiblc2 = 4.0342223672295e-08 wpdiblc2 = 3.61334755508028e-07 ppdiblc2 = -1.69607716833681e-13
+ pdiblcb = -1.29534565303 lpdiblcb = 6.77735757619769e-07 wpdiblcb = 6.26331982977302e-06 ppdiblcb = -3.34151244578305e-12
+ drout = 6.97636164512442 ldrout = -2.88716435586553e-06 wdrout = -2.63963994102197e-05 pdrout = 1.23114898409227e-11
+ pscbe1 = 913272503.407763 lpscbe1 = -290.478120948407 wpscbe1 = -1101.9889786158 ppscbe1 = 0.000636692282646369
+ pscbe2 = 2.51726455029538e-08 lpscbe2 = -4.69761650931152e-15 wpscbe2 = -4.74006211669815e-14 ppscbe2 = 2.08111901257703e-20
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.000338229425996697 lalpha0 = -9.95153693752968e-11 walpha0 = -7.21620346250065e-10 palpha0 = 1.7477830970355e-16
+ alpha1 = 6.35172826514999e-10 lalpha1 = -3.38867878809885e-16 walpha1 = -3.13165991488651e-15 palpha1 = 1.67075622289153e-21
+ beta0 = -181.540109506915 lbeta0 = 0.000130797633655794 wbeta0 = 0.00120282039956745 pbeta0 = -6.7028910184344e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -2.64426168013045e-08 lagidl = 1.35426873579305e-14 wagidl = 5.32436499156818e-14 pagidl = -8.46906329383715e-21
+ bgidl = -1790889707.00977 lbgidl = 1788.00086717409 wbgidl = 18003.6263811518 pbgidl = -0.00921923283791545
+ cgidl = -433.764839446938 lcgidl = 0.000127430853979789 wcgidl = -0.000360874463152782 pcgidl = 1.31020702999154e-9
+ egidl = 11.8225814421028 legidl = -5.67485391603844e-06 wegidl = -5.25314107930547e-05 pegidl = 2.69241815640172e-11
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.59725997543185 lkt1 = 9.78472520867404e-09 wkt1 = -8.52697815011454e-07 pkt1 = 3.5085880680722e-13
+ kt2 = -0.019032
+ at = 18000.0
+ ute = -0.795613480530498 lute = -3.13557122774126e-07 wute = -4.28787925922501e-06 pute = 2.17198308975899e-12
+ ua1 = 5.52e-10
+ ub1 = -5.05576226e-18 lub1 = 9.37134748521299e-25
+ uc1 = -4.1496e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 1.81e-6
+ sbref = 1.81e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.48 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 1.5e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.044948866372+0*(0.0/sqrt(l*w*mult))} wvth0 = 7.09593897057074e-8
+ k1 = 0.60838880728 wk1 = -3.8619255926156e-8
+ k2 = 0.027310130953636 wk2 = -2.03460883120647e-10
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 218738.3186 wvsat = -0.0549108812553517
+ ua = 2.726515265982e-09 wua = -5.39202498352478e-17
+ ub = -7.333429212e-19 wub = 5.87672179542007e-25
+ uc = -5.55395853e-11 wuc = 4.56193453686318e-17
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0192790399352 wu0 = -1.7828571114969e-10
+ a0 = 0.847939532084 wa0 = 1.77109249011854e-7
+ keta = -0.0063097319408 wketa = -4.73602857768804e-9
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.10342984253936 wags = 6.93614132000042e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.087664747963824+0*(0.009/sqrt(l*w*mult))} wvoff = -1.62341826790644e-8
+ nfactor = {1.87862710368+0*(0.02/sqrt(l*w*mult))} wnfactor = -4.13354582966494e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.476802e-05 wcit = -1.397223441612e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.63945410270796 wpclm = 2.11864061548752e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0045149854538708 wpdiblc2 = -4.61303854312952e-9
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 443756900.68032 wpscbe1 = -322.473804986034
+ pscbe2 = 1.501602017518e-08 wpscbe2 = -4.41382885205169e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 7.9767690028548e-05 walpha0 = -8.52762828170632e-11
+ alpha1 = 0.0
+ beta0 = 39.025870038368 wbeta0 = -2.22659292097783e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.95191799e-08 wagidl = -1.39023732440394e-14
+ bgidl = 1759488732.0 wbgidl = 47.5055970148078
+ cgidl = 1507.317328 wcgidl = -0.00148664574187517
+ egidl = 0.50431434165272 wegidl = 5.5441496418432e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.55692792 wkt1 = -5.58889376644797e-8
+ kt2 = -0.019032
+ at = 551054.95692 wat = -0.29964853928811
+ ute = -1.51702792 wute = -5.58889376644802e-8
+ ua1 = 2.2096e-11
+ ub1 = -3.5760173964e-18 wub1 = -2.54015221685063e-25
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.49 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 1.5e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.044948866372+0*(0.0/sqrt(l*w*mult))} wvth0 = 7.0959389705707e-8
+ k1 = 0.60838880728 wk1 = -3.86192559261564e-8
+ k2 = 0.027310130953636 wk2 = -2.03460883120647e-10
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 218738.3186 wvsat = -0.0549108812553515
+ ua = 2.726515265982e-09 wua = -5.39202498352494e-17
+ ub = -7.333429212e-19 wub = 5.87672179542007e-25
+ uc = -5.55395853e-11 wuc = 4.56193453686318e-17
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0192790399352 wu0 = -1.78285711149703e-10
+ a0 = 0.847939532084 wa0 = 1.77109249011853e-7
+ keta = -0.0063097319408 wketa = -4.73602857768804e-9
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.10342984253936 wags = 6.93614132000043e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.087664747963824+0*(0.009/sqrt(l*w*mult))} wvoff = -1.62341826790644e-8
+ nfactor = {1.87862710368+0*(0.02/sqrt(l*w*mult))} wnfactor = -4.13354582966493e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.476802e-05 wcit = -1.397223441612e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.63945410270796 wpclm = 2.11864061548752e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0045149854538708 wpdiblc2 = -4.61303854312952e-9
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 443756900.68032 wpscbe1 = -322.473804986034
+ pscbe2 = 1.501602017518e-08 wpscbe2 = -4.41382885205169e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 7.9767690028548e-05 walpha0 = -8.52762828170633e-11
+ alpha1 = 0.0
+ beta0 = 39.025870038368 wbeta0 = -2.22659292097781e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.95191799e-08 wagidl = -1.39023732440394e-14
+ bgidl = 1759488732.0 wbgidl = 47.5055970148078
+ cgidl = 1507.317328 wcgidl = -0.00148664574187517
+ egidl = 0.50431434165272 wegidl = 5.54414964184319e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.55692792 wkt1 = -5.58889376644802e-8
+ kt2 = -0.019032
+ at = 551054.95692 wat = -0.29964853928811
+ ute = -1.51702792 wute = -5.58889376644802e-8
+ ua1 = 2.2096e-11
+ ub1 = -3.5760173964e-18 wub1 = -2.54015221685063e-25
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.50 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 1.5e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.05587624115907+0*(0.0/sqrt(l*w*mult))} lvth0 = 8.66923825101163e-08 wvth0 = 8.65899721653847e-08 pvth0 = -1.24005304096764e-13
+ k1 = 0.625967126425871 lk1 = -1.39457682835361e-07 wk1 = -6.37633891023243e-08 pk1 = 1.99481106273798e-13
+ k2 = 0.0248597324759794 lk2 = 1.94402485744812e-08 wk2 = 3.30160380171025e-09 pk2 = -2.78074482024294e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 362995.80326267 lvsat = -1.14446747585872 wvsat = -0.261257652861743 pvsat = 1.63705314427317e-6
+ ua = 2.23520374332102e-09 lua = 3.8978224215885e-15 wua = 6.48854700048152e-16 pua = -5.57546857877472e-21
+ ub = -1.55621376550136e-19 lub = -4.58335676308742e-24 wub = -2.38704184254426e-25 pub = 6.55606101406082e-30
+ uc = -7.83491353785709e-11 luc = 1.80959679596092e-16 wuc = 7.824626265832e-17 puc = -2.58845811452328e-22
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0178672031329814 lu0 = 1.12008143295855e-08 wu0 = 1.84121412176463e-09 pu0 = -1.6021712021925e-14
+ a0 = 0.894725333139206 la0 = -3.71175386600481e-07 wa0 = 1.10186558467682e-07 pa0 = 5.30931500045649e-13
+ keta = -0.000473153646038265 lketa = -4.63045230843837e-08 wketa = -1.3084705189985e-08 pketa = 6.62342676470411e-14
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.0764637404057065 lags = 2.13935706107851e-07 wags = 1.07933887488595e-07 pags = -3.06014917630906e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0907545169764465+0*(0.009/sqrt(l*w*mult))} lvoff = 2.45126979104854e-08 wvoff = -1.18145585447951e-08 pvoff = -3.50631101673457e-14
+ nfactor = {1.90458153992707+0*(0.02/sqrt(l*w*mult))} lnfactor = -2.05909649738336e-07 wnfactor = -4.50479964300923e-07 pnfactor = 2.94534398443608e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.476802e-05 wcit = -1.397223441612e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -2.07807108031412 lpclm = 1.14132749849234e-05 wpclm = 4.17644697195725e-06 ppclm = -1.63256170180843e-11
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00768635955580281 lpdiblc2 = -2.51601122945482e-08 wpdiblc2 = -9.14939108677768e-09 ppdiblc2 = 3.59891755867955e-14
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 892749109.885198 lpscbe1 = -3562.08193668795 wpscbe1 = -964.714954985947 ppscbe1 = 0.00509522337473006
+ pscbe2 = -4.45815168992357e-08 lpscbe2 = 4.72817358367563e-13 wpscbe2 = 8.52045363279462e-14 ppscbe2 = -6.76320786313112e-19
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.000133797679699628 lalpha0 = -4.28647193205463e-10 walpha0 = -1.62561104222514e-10 palpha0 = 6.13139517044253e-16
+ alpha1 = 0.0
+ beta0 = 40.7443899152849 lbeta0 = -1.36338860361197e-05 wbeta0 = -4.68477406403902e-06 pbeta0 = 1.95019923893819e-11
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 2.98452416933394e-08 lagidl = -8.19218628677669e-14 wagidl = -2.86728339896028e-14 pagidl = 1.17181524177231e-19
+ bgidl = 1594079630.52902 lbgidl = 1312.27393356553 wbgidl = 284.107768213509 pbgidl = -0.00187708450821573
+ cgidl = 2160.5007716717 lcgidl = -0.00518203411628665 wcgidl = -0.00242096325880383 pcgidl = 7.41241269214113e-9
+ egidl = 1.51825613067546 legidl = -8.04411225292086e-06 wegidl = -8.95933454484542e-07 pegidl = 1.15063464312515e-11
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.55692792 wkt1 = -5.58889376644802e-8
+ kt2 = -0.019032
+ at = 972050.897644166 lat = -3.33997340071487 wat = -0.901843658875601 pat = 4.77751799222296e-6
+ ute = -1.4786053644899 lute = -3.04825536252154e-07 wute = -1.1084879160146e-07 pute = 4.36024276008301e-13
+ ua1 = 2.2096e-11
+ ub1 = -3.40138688160659e-18 lub1 = -1.38543206226606e-24 wub1 = -5.03807757828635e-25 pub1 = 1.98173033445773e-30
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.51 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 1.5e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.0066965220918+0*(0.0/sqrt(l*w*mult))} lvth0 = -1.0675628833959e-07 wvth0 = 2.15033629183089e-08 pvth0 = 1.32013198809656e-13
+ k1 = 0.623224775543493 lk1 = -1.28670631927775e-07 wk1 = -5.9840713946066e-08 pk1 = 1.84051243933281e-13
+ k2 = 0.0267815550317242 lk2 = 1.1880749942346e-08 wk2 = 3.51232809535252e-09 pk2 = -2.86363332650927e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 50700.431713587 lvsat = 0.0839479296064581 wvsat = 0.185451520374295 pvsat = -1.20079622196655e-7
+ ua = 3.84197097774937e-09 lua = -2.42240452887159e-15 wua = -1.67954206928073e-15 pua = 3.5832917553643e-21
+ ub = -3.38336767530554e-18 lub = 8.11299944179848e-24 wub = 4.27946512868534e-24 pub = -1.12161805692343e-29
+ uc = -9.73356634674913e-11 luc = 2.55643282766501e-16 wuc = 1.23287704147372e-16 puc = -4.36016546756723e-22
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0189415386347081 lu0 = 6.97491026186602e-09 wu0 = 1.27058701714887e-10 pu0 = -9.27907310638222e-15
+ a0 = 0.574457872731588 la0 = 8.88598270250187e-07 wa0 = 7.05487314169824e-07 pa0 = -1.81068699901251e-12
+ keta = -0.000618437305182441 lketa = -4.57330490847218e-08 wketa = -1.28768905722432e-08 pketa = 6.54168278090806e-14
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.0511632542832482 lags = 3.13455294772971e-07 wags = 1.23680595681081e-07 pags = -3.67954673039592e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0300976774548448+0*(0.009/sqrt(l*w*mult))} lvoff = -2.14081283631933e-07 wvoff = -9.85784657375313e-08 pvoff = 3.06223152594818e-13
+ nfactor = {2.75610578772633+0*(0.02/sqrt(l*w*mult))} lnfactor = -3.55538453607796e-06 wnfactor = -1.571318759541e-06 pnfactor = 4.70335940371441e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.476802e-05 wcit = -1.397223441612e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -0.040495968954438 leta0 = 4.73971496362127e-07 weta0 = 1.72358156968242e-07 peta0 = -6.77971672225364e-13
+ etab = -0.173671860938041 letab = 4.07793783359089e-07 wetab = 1.48292851916939e-07 petab = -5.8331067447954e-13
+ dsub = 1.06398666638702 ldsub = -1.98243407216667e-06 wdsub = -7.20905551519989e-07 pdsub = 2.83568559143164e-12
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.25160391944343 lpclm = -1.68401827499793e-06 wpclm = -5.86340125745954e-07 ppclm = 2.40882984466669e-12
+ pdiblc1 = 0.768990796247144 lpdiblc1 = -1.49076219199212e-06 wpdiblc1 = -5.42110708896692e-07 ppdiblc1 = 2.13239518399868e-12
+ pdiblc2 = -0.00350439484448231 lpdiblc2 = 1.88587760927454e-08 wpdiblc2 = 6.85793115191656e-09 ppdiblc2 = -2.69757064757196e-14
+ pdiblcb = 0.352730310202 lpdiblcb = -1.48580406383112e-06 wpdiblcb = -5.40307702094802e-07 ppdiblcb = 2.12530304772841e-12
+ drout = -0.2710066824444 ldrout = 3.26876894042846e-06 wdrout = 1.18867694460856e-06 pdrout = -4.67566670500251e-12
+ pscbe1 = -519638603.384229 lpscbe1 = 1993.55219539591 wpscbe1 = 1055.57290440092 ppscbe1 = -0.00285158902160748
+ pscbe2 = 1.35075743556534e-07 lpscbe2 = -2.3386537392151e-13 wpscbe2 = -1.7177828697155e-13 ppscbe2 = 3.34522434049571e-19
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 6.74001869113994e-05 lalpha0 = -1.67472323335501e-10 walpha0 = -6.75857321532751e-11 palpha0 = 2.39553416133041e-16
+ alpha1 = -1.88865155101e-10 lalpha1 = 7.42902031915559e-16 walpha1 = 2.70153851047401e-16 palpha1 = -1.06265152386421e-21
+ beta0 = 102.194102760424 lbeta0 = -0.000255346638761039 wbeta0 = -9.25828120160033e-05 pbeta0 = 3.65249364163623e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.85841638885338e-08 lagidl = -3.7626357017175e-14 wagidl = -2.6669976211595e-14 pagidl = 1.09303273093148e-19
+ bgidl = 2962729308.7943 lbgidl = -4071.31641913933 wbgidl = -1408.24830164199 pbgidl = 0.0047798065543412
+ cgidl = 1879.50441278018 lcgidl = -0.00407673353360508 wcgidl = -0.00303126953907623 pcgidl = 9.81305549712402e-9
+ egidl = -3.99107690641203 legidl = 1.3626876795128e-05 wegidl = 6.98464957776362e-06 pegidl = -1.94919663290118e-11
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.55328517724495 lkt1 = -1.43287468407038e-08 wkt1 = -6.93966302168497e-08 pkt1 = 5.31325761932101e-14
+ kt2 = -0.019032
+ at = 186192.275225939 lat = -0.248794580139664 wat = 0.291492458009272 pat = 8.35244097757264e-8
+ ute = -1.6219898287096 lute = 2.59177970678354e-07 wute = -1.0806154041896e-07 pute = 4.25060609545684e-13
+ ua1 = -4.9057671776e-10 lua1 = 2.01660069867255e-15 pua1 = -9.4039548065783e-38
+ ub1 = -3.51850269508741e-18 lub1 = -9.24756424360198e-25 wub1 = 3.54171698723141e-25 pub1 = -1.39313614778597e-30
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.52 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 1.5e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.12298031258001+0*(0.0/sqrt(l*w*mult))} lvth0 = 1.18079001988319e-07 wvth0 = 1.67538036609499e-07 pvth0 = -1.50345572945631e-13
+ k1 = 0.537254513963487 lk1 = 3.75532986884748e-08 wk1 = 6.31316640395441e-08 pk1 = -5.37164637637864e-14
+ k2 = 0.0250423688449188 lk2 = 1.52434751304653e-08 wk2 = -2.22237780142922e-09 pk2 = -1.75482507401357e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 228483.024768909 lvsat = -0.259795602978971 wvsat = -0.0287910328366953 pvsat = 2.9415942564956e-7
+ ua = 4.33395301289895e-09 lua = -3.37365425374349e-15 wua = -2.29914853390855e-15 pua = 4.7813039527545e-21
+ ub = 5.69536393456433e-19 lub = 4.70039660326849e-25 wub = -1.27797687115243e-24 pub = -4.70838675337982e-31
+ uc = 6.72094616399826e-11 luc = -6.25055393544249e-17 wuc = -1.95349455332172e-16 puc = 1.80069994282773e-22
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0297758696252904 lu0 = -1.39733228800798e-08 wu0 = -1.45775261030279e-08 pu0 = 1.91523151365119e-14
+ a0 = 1.21968214625285 la0 = -3.58946088724533e-07 wa0 = -4.76945188120721e-07 pa0 = 4.75552156328769e-13
+ keta = 0.0989231592624551 lketa = -2.38197223756232e-07 wketa = -1.55261787552171e-07 pketa = 3.40718738044256e-13
+ a1 = 0.0
+ a2 = 0.5
+ ags = -0.654301490283014 lags = 1.67747490571556e-06 wags = 1.1553486215677e-06 pags = -2.3626899594315e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.218613910572313+0*(0.009/sqrt(l*w*mult))} lvoff = 1.50415795681857e-07 wvoff = 1.71076285211094e-07 pvoff = -2.15155656638103e-13
+ nfactor = {0.0736966582119569+0*(0.02/sqrt(l*w*mult))} lnfactor = 1.63106692788373e-06 wnfactor = 2.21132344488062e-06 pnfactor = -2.61039821174581e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 2.38865155101e-05 lcit = -1.76306566612559e-11 wcit = -2.70153851047401e-11 pcit = 2.52189970722004e-17
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.450885088820161 leta0 = -4.76116235750349e-07 weta0 = -5.30516256358891e-07 peta0 = 6.81039520314714e-13
+ etab = 0.00968478473468184 letab = 5.32727921676508e-08 wetab = -1.13981594193197e-07 petab = -7.62017215533608e-14
+ dsub = 0.028031281693754 ldsub = 2.05908439146808e-08 wdsub = 7.60931246477564e-07 pdsub = -2.94532666806228e-14
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.708883550884292 lpclm = 2.10659405131806e-06 wpclm = 2.21795590578782e-06 ppclm = -3.01329055378402e-12
+ pdiblc1 = -0.385354879619772 lpdiblc1 = 7.41170944024938e-07 wpdiblc1 = 1.1090722719374e-06 ppdiblc1 = -1.06017536535894e-12
+ pdiblc2 = 0.0104845338457042 lpdiblc2 = -8.1888874743736e-09 wpdiblc2 = -1.31519163800983e-08 ppdiblc2 = 1.17134337766689e-14
+ pdiblcb = -0.780460620404 lpdiblcb = 7.05226266450236e-07 wpdiblcb = 1.0806154041896e-06 ppdiblcb = -1.00875988288802e-12
+ drout = 2.49431095379388 ldrout = -2.07798653582643e-06 wdrout = -2.76684999417248e-06 pdrout = 2.97236440876534e-12
+ pscbe1 = 637008906.210778 lpscbe1 = -242.831547643583 wpscbe1 = -598.902633208834 ppscbe1 = 0.000347347702738667
+ pscbe2 = 1.41008009285865e-08 lpscbe2 = 4.02825243396361e-17 wpscbe2 = 1.26499681312226e-15 ppscbe2 = -5.762036451056e-23
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -0.000142886356161136 lalpha0 = 2.39117759127961e-10 walpha0 = 2.33209400776937e-10 palpha0 = -3.4203547736319e-16
+ alpha1 = 3.77730310202e-10 lalpha1 = -3.52613133225118e-16 walpha1 = -5.40307702094802e-16 palpha1 = 5.04379941444008e-22
+ beta0 = -115.862765471532 lbeta0 = 0.00016626740624979 wbeta0 = 0.000219327040644197 pbeta0 = -2.37829895504137e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -1.8018710524206e-09 lagidl = 1.79014347133499e-15 wagidl = 4.16007981582428e-14 pagidl = -2.26986105048047e-20
+ bgidl = 214501140.229973 lbgidl = 1242.39648592063 wbgidl = 2006.60486021684 pbgidl = -0.00182282910837865
+ cgidl = -1607.75372506741 lcgidl = 0.00266589751221393 wcgidl = 0.00484944945434949 pcgidl = -5.42435408025959e-9
+ egidl = 5.28345645987543 legidl = -4.30547984125566e-06 wegidl = -6.28169859657415e-06 pegidl = 6.15858419781114e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.4692944304091 lkt1 = -1.76725275801553e-07 wkt1 = -1.59305059445941e-07 pkt1 = 2.26970973649804e-13
+ kt2 = -0.019032
+ at = 65400.0829306645 lat = -0.0152422723757899 wat = 0.699299137553425 pat = -7.0497184415629e-7
+ ute = -1.4509697819394 lute = -7.14901448520608e-08 wute = 3.35189711972385e-08 pute = 1.51313982433202e-13
+ ua1 = 5.524e-10
+ ub1 = -4.37567587332518e-18 lub1 = 7.3259220162842e-25 wub1 = -7.08343397446285e-25 pub1 = 6.61242103233096e-31
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.81e-6
+ sbref = 2.81e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.53 pmos
* DC IV MOS Parameters
+ lmin = 8.0e-07 lmax = 1e-06 wmin = 1.5e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.866660657676803+0*(0.0/sqrt(l*w*mult))} lvth0 = -1.21196677462101e-07 wvth0 = -2.67690207432878e-07 pvth0 = 2.55942169009148e-13
+ k1 = 0.583914026381164 lk1 = -6.00358945098726e-09 wk1 = 1.962961797984e-08 pk1 = -1.31070862568235e-14
+ k2 = 0.0324290626975307 lk2 = 8.34795948558284e-09 wk2 = -3.53177847696432e-08 pk2 = 1.33464771417269e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -443542.08696275 lvsat = 0.367543198948091 wvsat = 1.33781772020582 pvsat = -9.81576678359389e-7
+ ua = -8.77907755197037e-09 lua = 8.86742534371486e-15 wua = 2.29661165799134e-14 pua = -1.88039473573239e-20
+ ub = 1.01963127998152e-17 lub = -8.51660424889114e-24 wub = -2.03976897550272e-23 pub = 1.73775089003235e-29
+ uc = 1.22316471485258e-11 luc = -1.11834746375775e-17 wuc = -1.73506795375307e-17 puc = 1.39072470845967e-23
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = -0.00855746916733047 lu0 = 2.18110405495257e-08 wu0 = 5.59957570872317e-08 pu0 = -4.67281975880113e-14
+ a0 = 0.638447544086397 la0 = 1.83639318570857e-07 wa0 = 6.38420623216997e-07 pa0 = -5.65647405384047e-13
+ keta = -0.488169854084381 lketa = 3.09857039668107e-07 wketa = 9.73032907996342e-07 pketa = -7.12550001723759e-13
+ a1 = 0.0
+ a2 = 0.5
+ ags = 2.73979819579286 lags = -1.4909341217347e-06 wags = -6.57062730196477e-06 pags = 4.84954719506568e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0389825658247304+0*(0.009/sqrt(l*w*mult))} lvoff = -1.72709627967346e-08 wvoff = -1.66653488112407e-07 pvoff = 1.00116775408252e-13
+ nfactor = {1.8635265758288+0*(0.02/sqrt(l*w*mult))} lnfactor = -3.97482493611806e-08 wnfactor = -8.3951326789854e-07 pnfactor = 2.37573113817104e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -1.3337625e-05 lcit = 1.7118264625625e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -0.257295347870041 leta0 = 1.84973742802138e-07 weta0 = 8.66353177770058e-07 peta0 = -6.22945080791831e-13
+ etab = 0.301059117623448 letab = -2.18726604455677e-07 wetab = -8.7650872100038e-07 petab = 6.35621163956778e-13
+ dsub = -0.807767752762231 ldsub = 8.00813421574515e-07 wdsub = 3.5029681389142e-06 pdsub = -2.58915841595468e-12
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 4.28982414943843 lpclm = -2.55972458047169e-06 wpclm = -6.56370603867539e-06 ppclm = 5.18443477968211e-12
+ pdiblc1 = 0.221424537533376 lpdiblc1 = 1.7473932421539e-07 wpdiblc1 = -9.53185928311056e-08 ppdiblc1 = 6.41295288567871e-14
+ pdiblc2 = -0.0506705204649743 lpdiblc2 = 4.88996614999163e-08 wpdiblc2 = 4.64493346005113e-08 ppdiblc2 = -4.39246320199851e-14
+ pdiblcb = -0.025
+ drout = 0.0684654035908228 ldrout = 1.86552414515872e-07 wdrout = 7.7602262624747e-07 pdrout = -3.34924896759791e-13
+ pscbe1 = 183388895.767649 lpscbe1 = 180.625000205131 wpscbe1 = -740.12417018079 ppscbe1 = 0.000479178713609673
+ pscbe2 = 1.64250625835055e-08 lpscbe2 = -2.12942735183552e-15 wpscbe2 = 5.81365146809237e-15 ppscbe2 = -4.30381222819843e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.00051864859907065 lalpha0 = -3.78428429255687e-10 walpha0 = -7.77605892697802e-10 palpha0 = 6.01565653171947e-16
+ alpha1 = 0.0
+ beta0 = 131.581937267725 lbeta0 = -6.4723460980821e-05 wbeta0 = -0.000186966267496339 pbeta0 = 1.41446939111593e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -9.20334616358777e-08 lagidl = 8.60217844389451e-14 wagidl = 1.72413810920868e-13 pagidl = -1.44813211983779e-19
+ bgidl = 519453177.916199 lbgidl = 957.722233980352 wbgidl = 443.383569451275 pbgidl = -0.000363554217342538
+ cgidl = 3883.1701903734 lcgidl = -0.00245990741746964 wcgidl = -0.00438435679883136 pcgidl = 3.195450226116e-9
+ egidl = 0.253669756486135 legidl = 3.89851195291764e-07 wegidl = 4.74145502936085e-06 pegidl = -4.13158482776731e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.725020102803001 lkt1 = 6.19959180065156e-08 wkt1 = 3.91294520658602e-07 pkt1 = -2.87016487375689e-13
+ kt2 = -0.019032
+ at = 119870.2026515 lat = -0.0660904014857886 wat = -0.209619494745422 pat = 1.43508243687844e-7
+ ute = -1.702684960707 lute = 1.63487233103388e-07 wute = 9.13020548203407e-07 pute = -6.69705137209942e-13
+ ua1 = 5.524e-10
+ ub1 = -3.5909e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.41e-6
+ sbref = 2.41e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.54 pmos
* DC IV MOS Parameters
+ lmin = 6e-07 lmax = 8.0e-07 wmin = 1.5e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.04643154363682+0*(0.0/sqrt(l*w*mult))} lvth0 = 1.06661662440006e-08 wvth0 = 6.19187258468181e-08 pvth0 = 1.4172368403825e-14
+ k1 = 0.703909422363938 lk1 = -9.40208123813338e-08 wk1 = -3.73859504771822e-07 pk1 = 2.75519152727134e-13
+ k2 = 0.00700690189381281 lk2 = 2.69952415459139e-08 wk2 = 7.60298264724776e-08 pk2 = -6.83275524424249e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 19846.0998206937 lvsat = 0.0276456470015007 wvsat = -0.0158326626233596 pvsat = 1.13326456977252e-8
+ ua = 2.86014021186557e-09 lua = 3.30000917852369e-16 wua = -1.26942333753074e-15 pua = -1.02705765017899e-21
+ ub = -1.43399870057557e-19 lub = -9.32373306976082e-25 wub = 1.18813618979497e-24 pub = 1.54419764066675e-30
+ uc = -5.21290375615217e-12 luc = 1.61219067375828e-18 wuc = 8.05012932965085e-18 puc = -4.72437322352529e-24
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0248513743929271 lu0 = -2.69451324614096e-09 wu0 = -9.42706030099514e-09 pu0 = 1.25976608034e-15
+ a0 = 1.0058192654646 la0 = -8.58296759186617e-08 wa0 = -4.75632045373058e-07 pa0 = 2.51515797290102e-13
+ keta = -0.147837369708223 lketa = 6.02214607157729e-08 wketa = 6.89280665851459e-08 pketa = -4.9384580024439e-14
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.672752152126146 lags = 2.52544865250561e-08 wags = 1.41737431616628e-07 pags = -7.40058988399447e-14
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0532502144231446+0*(0.009/sqrt(l*w*mult))} lvoff = -6.8055712115546e-09 wvoff = -5.73513174435164e-08 pvoff = 1.99430867117669e-14
+ nfactor = {2.21462896624637+0*(0.02/sqrt(l*w*mult))} lnfactor = -2.9728360824442e-07 wnfactor = -1.64068183874832e-06 pnfactor = 8.25234266378269e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.0254482126818668 leta0 = -2.24200725804892e-08 weta0 = -6.88172625354335e-08 peta0 = 6.30071130244488e-14
+ etab = 0.0105088180835521 letab = -5.60650699166545e-09 wetab = -3.65118272030281e-08 petab = 1.94792423719515e-14
+ dsub = 0.300836798761218 ldsub = -1.23535599906928e-08 wdsub = -7.62020600368663e-08 pdsub = 3.61808208269175e-14
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.665762758130082 lpclm = 9.85425703599319e-08 wpclm = 8.97989580016482e-07 ppclm = -2.88756265106471e-13
+ pdiblc1 = 0.318271163185807 lpdiblc1 = 1.03701840066203e-07 wpdiblc1 = 4.06406716741192e-07 ppdiblc1 = -3.03888494341042e-13
+ pdiblc2 = 0.0191607476168585 lpdiblc2 = -2.32192279444851e-09 wpdiblc2 = -2.27101237649719e-08 ppdiblc2 = 6.80417648838867e-15
+ pdiblcb = -0.025
+ drout = 0.567475791143008 ldrout = -1.79474199805593e-07 wdrout = -3.97598778808116e-07 pdrout = 5.25932271955508e-13
+ pscbe1 = 352309139.173831 lpscbe1 = 56.7211570654792 wpscbe1 = 139.753584710172 ppscbe1 = -0.000166216018991622
+ pscbe2 = 1.63987542339712e-08 lpscbe2 = -2.11013004591037e-15 wpscbe2 = -8.48393338206472e-15 ppscbe2 = 6.18353774731603e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -4.39313461157129e-06 lalpha0 = 5.22529760889048e-12 walpha0 = 6.33943685639822e-11 palpha0 = -1.53122434648783e-17
+ alpha1 = 0.0
+ beta0 = 45.1938441508515 lbeta0 = -1.35736273912827e-06 wbeta0 = 4.48017609659993e-07 pbeta0 = 3.9776239149179e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.51189942640194e-07 lagidl = -9.23837987145748e-14 wagidl = -3.54914092915548e-13 pagidl = 2.41984442119751e-19
+ bgidl = 1215138144.87802 lbgidl = 447.433832289023 wbgidl = 1735.27465322058 pbgidl = -0.00131116278674274
+ cgidl = 1689.4917446056 lcgidl = -0.000850833309106732 wcgidl = -0.00342708562534272 pcgidl = 2.49328703400622e-9
+ egidl = 3.4588638211966 legidl = -1.96117467714368e-06 wegidl = -8.72624167170762e-06 pegidl = 5.74703804094991e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.647565825580799 lkt1 = 5.18281839264435e-09 wkt1 = 5.96340553773758e-08 pkt1 = -4.3741877789582e-14
+ kt2 = -0.019032
+ at = 40809.4074697 lat = -0.00809891291596231 wat = 0.00839053635039633 pat = -1.64032041710936e-8
+ ute = -1.24448848507739 lute = -1.7260217275331e-07 wute = -8.65439228664183e-07 pute = 6.3480400142132e-13
+ ua1 = 5.5346701e-10 lua1 = -7.8265717005015e-19
+ ub1 = -7.32454158061033e-19 lub1 = -2.09668431729144e-24 wub1 = -1.06566056959372e-23 pub1 = 7.81667356099845e-30
+ uc1 = -4.62025009583811e-10 luc1 = 2.58798908654773e-16 wuc1 = 5.0468301065874e-16 puc1 = -3.70187511733239e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.02e-6
+ sbref = 2.01e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.55 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 6e-07 wmin = 1.5e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.014/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.746647037564705+0*(0.0/sqrt(l*w*mult))} lvth0 = -1.49270366668005e-07 wvth0 = -1.32986006072795e-07 pvth0 = 1.18155017406597e-13
+ k1 = 0.440035016470969 lk1 = 4.67575025345959e-08 wk1 = 4.95818872568352e-07 pk1 = -1.88458609975735e-13
+ k2 = 0.121914379697615 lk2 = -3.43084723998037e-08 wk2 = -2.4604215237391e-07 pk2 = 1.03499458632017e-13
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -436710.994284636 lvsat = 0.271221139492165 wvsat = 0.695453115884577 pvsat = -3.68141873565152e-7
+ ua = 3.51719082209898e-09 lua = -2.0538867960208e-17 wua = -6.79342135214238e-15 pua = 1.92002291060639e-21
+ ub = -1.07694867609421e-17 lub = 4.73669717974525e-24 wub = 2.02338971757677e-23 pub = -8.61681107415461e-30
+ uc = 2.78023097920593e-10 luc = -1.49495632400794e-16 wuc = -3.95946097421507e-16 puc = 2.10809633729351e-22
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0038315093420381 lu0 = 8.51968985783354e-09 wu0 = 6.78861487652279e-09 pu0 = -7.3913777052417e-15
+ a0 = 0.0385705972920363 la0 = 4.30202324794741e-07 wa0 = 1.31393995571465e-06 pa0 = -7.03229813150197e-13
+ keta = -0.37777374642199 lketa = 1.82893667374451e-07 wketa = 4.45829840263382e-07 pketa = -2.50463560790646e-13
+ a1 = 0.0
+ a2 = 0.5
+ ags = 5.73122677842882 lags = -2.67346701898055e-06 wags = -7.93458713177556e-06 pags = 4.23475363735261e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {0.288681625762145+0*(0.009/sqrt(l*w*mult))} lvoff = -1.89227917609608e-07 wvoff = -4.54768686338037e-07 pvoff = 2.31967240103839e-13
+ nfactor = {4.73460357597905+0*(0.02/sqrt(l*w*mult))} lnfactor = -1.64170266240985e-06 wnfactor = -4.5317206472773e-06 pnfactor = 2.36761792592253e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -1.06116696023258 leta0 = 5.57294555245233e-07 weta0 = 1.28667527857213e-06 peta0 = -6.60154935119142e-13
+ etab = 0.0702190071260886 letab = -3.74621913968039e-08 wetab = -1.38463785365604e-08 petab = 7.38711218114764e-15
+ dsub = 0.129929717509807 ldsub = 7.88262223923419e-08 wdsub = 1.91732994950558e-07 pdsub = -1.06763870684148e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 3.68634050504328 lpclm = -1.51295076050699e-06 wpclm = -3.2974334292763e-06 ppclm = 1.94952288746628e-12
+ pdiblc1 = 1.90456671834687 lpdiblc1 = -7.42594770089998e-07 wpdiblc1 = -8.42324425956965e-07 ppdiblc1 = 3.6231581394414e-13
+ pdiblc2 = 0.0626333303928824 lpdiblc2 = -2.55147630683712e-08 wpdiblc2 = -5.37797777788954e-08 ppdiblc2 = 2.33799922530869e-14
+ pdiblcb = 1.66879420404 lpdiblcb = -9.0364767682636e-07 wpdiblcb = -2.42281339222404e-06 ppdiblcb = 1.29258305881849e-12
+ drout = -3.10228027851842 ldrout = 1.77835901213913e-06 wdrout = 3.13811335467484e-06 pdrout = -1.36038782981832e-12
+ pscbe1 = 737294099.809321 lpscbe1 = -148.670244358358 wpscbe1 = -586.300808840505 ppscbe1 = 0.000221137630239631
+ pscbe2 = 4.19896300065785e-09 lpscbe2 = 4.39851957601848e-15 wpscbe2 = 1.40607838798414e-14 ppscbe2 = -5.84418163549722e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.00010400882762687 lalpha0 = -5.26076912551291e-11 walpha0 = -3.52588994635334e-11 palpha0 = 3.73197682941414e-17
+ alpha1 = -8.4689710202e-10 lalpha1 = 4.5182383841318e-16 walpha1 = 1.21140669611202e-15 palpha1 = -6.46291529409243e-22
+ beta0 = 392.140637703709 lbeta0 = -0.000186455211833546 wbeta0 = -0.000478297104143045 pbeta0 = 2.59390540095595e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -2.20252492233001e-07 lagidl = 1.05782597502449e-13 wagidl = 6.21185271739977e-13 pagidl = -2.78769449420795e-19
+ bgidl = 7598507694.1551 lbgidl = -2958.12573909805 wbgidl = -9511.1200996061 pbgidl = 0.00468884504586406
+ cgidl = -3935.57636025128 lcgidl = 0.00215016865017494 wcgidl = 0.00990085502828139 pcgidl = -4.61723594440551e-9
+ egidl = -15.4418823144363 legidl = 8.12246788994713e-06 wegidl = 2.73645373858899e-05 pegidl = -1.35075730401737e-11
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -1.0294351247272 lkt1 = 2.08911998833745e-07 wkt1 = 4.13750835534537e-07 pkt1 = -2.32664950587329e-13
+ kt2 = -0.019032
+ at = 4959.22689900003 lat = 0.011027337669409 wat = 0.0382147597398089 pat = -3.23145764704621e-8
+ ute = -2.96195505159466 lute = 7.43674827816488e-07 wute = 2.06038107867083e-06 pute = -9.26135761643448e-13
+ ua1 = 5.52e-10
+ ub1 = -9.29459000005112e-18 lub1 = 2.47125796508948e-24 wub1 = 1.24214862424122e-23 pub1 = -4.49560387857069e-30
+ uc1 = 2.3066805216e-11 wuc1 = -1.89195231781798e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 1.81e-6
+ sbref = 1.81e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.56 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 1e-06 wmax = 1.5e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.998223397788+0*(0.0/sqrt(l*w*mult))} wvth0 = 4.12299909034219e-9
+ k1 = 0.57495159048 wk1 = 9.20953960786497e-9
+ k2 = 0.02861232770688 wk2 = -2.0661309321414e-9
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 366792.197528 wvsat = -0.266688037997236
+ ua = 3.4926324127468e-09 wua = -1.1497788132705e-15
+ ub = -1.394212341656e-18 wub = 1.53298376377879e-24
+ uc = 1.6288969324584e-11 wuc = -5.71246501377009e-17
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.02093646243616 wu0 = -2.54907280105787e-9
+ a0 = 1.0844520545876 wa0 = -1.6119968225243e-7
+ keta = -0.0122980363056 wketa = 3.82967791554807e-9
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.16065182485016 wags = -1.2489253629258e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.082888250244452+0*(0.009/sqrt(l*w*mult))} wvoff = -2.30665136758404e-8
+ nfactor = {1.62506125236+0*(0.02/sqrt(l*w*mult))} wnfactor = -5.06524678432593e-8
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 5.0e-6
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.25248730812388 wpclm = -2.01800973021481e-6
+ pdiblc1 = 0.39
+ pdiblc2 = -0.0027071481060792 wpdiblc2 = 5.71754463382433e-9
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 206400231.27768 wpscbe1 = 17.0425990675187
+ pscbe2 = 1.495993038928e-08 wpscbe2 = 3.60928777695451e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -6.1895678072668e-05 walpha0 = 1.17359848895125e-10
+ alpha1 = 0.0
+ beta0 = 34.547362338112 wbeta0 = 4.17949136451458e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -9.1802824e-09 wagidl = 2.71495098266544e-14
+ bgidl = 2299399107.6 wbgidl = -724.785443705687
+ cgidl = -1266.276784 wcgidl = 0.0024807199174943
+ egidl = -0.27673521064156 wegidl = 1.67163293008337e-6
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.67043248 wkt1 = 1.0646866598688e-7
+ kt2 = -0.019032
+ at = 696017.46976 wat = -0.507003787429523
+ ute = -1.5561
+ ua1 = 2.2096e-11
+ ub1 = -5.0131836428e-18 wub1 = 1.80171600016298e-24
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.57 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 1e-06 wmax = 1.5e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.998223397788+0*(0.0/sqrt(l*w*mult))} wvth0 = 4.12299909034261e-9
+ k1 = 0.57495159048 wk1 = 9.2095396078654e-9
+ k2 = 0.02861232770688 wk2 = -2.06613093214138e-9
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 366792.197528 wvsat = -0.266688037997237
+ ua = 3.4926324127468e-09 wua = -1.1497788132705e-15
+ ub = -1.394212341656e-18 wub = 1.53298376377879e-24
+ uc = 1.6288969324584e-11 wuc = -5.71246501377009e-17
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.02093646243616 wu0 = -2.54907280105788e-9
+ a0 = 1.0844520545876 wa0 = -1.61199682252431e-7
+ keta = -0.0122980363056 wketa = 3.82967791554807e-9
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.16065182485016 wags = -1.2489253629258e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.082888250244452+0*(0.009/sqrt(l*w*mult))} wvoff = -2.30665136758404e-8
+ nfactor = {1.62506125236+0*(0.02/sqrt(l*w*mult))} wnfactor = -5.06524678432584e-8
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 5.0e-6
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.25248730812388 wpclm = -2.01800973021481e-6
+ pdiblc1 = 0.39
+ pdiblc2 = -0.0027071481060792 wpdiblc2 = 5.71754463382432e-9
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 206400231.27768 wpscbe1 = 17.0425990675188
+ pscbe2 = 1.495993038928e-08 wpscbe2 = 3.60928777695451e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -6.1895678072668e-05 walpha0 = 1.17359848895125e-10
+ alpha1 = 0.0
+ beta0 = 34.547362338112 wbeta0 = 4.17949136451455e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -9.1802824e-09 wagidl = 2.71495098266544e-14
+ bgidl = 2299399107.6 wbgidl = -724.785443705685
+ cgidl = -1266.276784 wcgidl = 0.0024807199174943
+ egidl = -0.27673521064156 wegidl = 1.67163293008337e-6
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.67043248 wkt1 = 1.0646866598688e-7
+ kt2 = -0.019032
+ at = 696017.46976 wat = -0.507003787429523
+ ute = -1.5561
+ ua1 = 2.2096e-11
+ ub1 = -5.0131836428e-18 wub1 = 1.80171600016298e-24
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.58 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 1e-06 wmax = 1.5e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.975682956561988+0*(0.0/sqrt(l*w*mult))} lvth0 = -1.78824703168773e-07 wvth0 = -2.81189832819931e-08 pvth0 = 2.55791928360829e-13
+ k1 = 0.612006626591929 lk1 = -2.93976314269168e-07 wk1 = -4.37942063768541e-08 pk1 = 4.20505483788502e-13
+ k2 = 0.0163668112238949 lk2 = 9.71498662453452e-08 wk2 = 1.54499293182195e-08 pk2 = -1.38963751576539e-13
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 440122.741584762 lvsat = -0.581768237927043 wvsat = -0.371580488199293 pvsat = 8.3216477814027e-7
+ ua = 2.99045066914882e-09 lua = 3.98406137374331e-15 wua = -4.31455034137487e-16 pua = -5.69882529337065e-21
+ ub = -1.20796366582665e-18 lub = -1.47760480093552e-24 wub = 1.26657254038044e-24 pub = 2.11357477288698e-30
+ uc = 4.41150506943009e-11 luc = -2.20758355677056e-16 wuc = -9.69272438854322e-17 puc = 3.15774076510595e-22
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0194044517036351 lu0 = 1.21542148065398e-08 wu0 = -3.57675457189892e-10 pu0 = -1.73854617845635e-14
+ a0 = 1.03015828372507 la0 = 4.30739902606727e-07 wa0 = -8.35375466480452e-08 pa0 = -6.16132941128077e-13
+ keta = -0.0153087351162151 lketa = 2.38853940675092e-08 wketa = 8.13619955844481e-09 pketa = -3.41658109865295e-14
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.172085471896507 lags = -9.07088960104286e-08 wags = -2.8844010966235e-08 pags = 1.29750549106693e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0634738834874204+0*(0.009/sqrt(l*w*mult))} lvoff = -1.54023975738744e-07 wvoff = -5.08369403712989e-08 pvoff = 2.20316819040553e-13
+ nfactor = {1.74389355088388+0*(0.02/sqrt(l*w*mult))} lnfactor = -9.42756634500733e-07 wnfactor = -2.20630900645614e-07 pnfactor = 1.34852474652964e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.4149391632575e-05 lcit = -7.2586744263992e-11 wcit = -1.30873446875851e-11 pcit = 1.0382851451568e-16
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 3.77145305764444 lpclm = -1.20507223686501e-05 wpclm = -4.19074745212352e-06 ppclm = 1.72374255804514e-11
+ pdiblc1 = 0.39
+ pdiblc2 = -0.00663784862132997 lpdiblc2 = 3.11842321912445e-08 wpdiblc2 = 1.13400422350421e-08 ppdiblc2 = -4.46061128317493e-14
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 207024329.579721 lpscbe1 = -4.9512869997352 wpscbe1 = 16.1498851116892 ppscbe1 = 7.08235063214338e-6
+ pscbe2 = 1.49757881148576e-08 lpscbe2 = -1.25807345158376e-16 wpscbe2 = 1.34098919570136e-17 ppscbe2 = 1.79955581358635e-22
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -0.000179451711488819 lalpha0 = 9.32631378887204e-10 walpha0 = 2.85512704429788e-10 palpha0 = -1.33404152014853e-15
+ alpha1 = 1.829878326515e-10 lalpha1 = -1.45173488527984e-15 walpha1 = -2.61746893751702e-16 palpha1 = 2.07657029031359e-21
+ beta0 = -31.4004973530022 lbeta0 = 0.000523197674598753 wbeta0 = 9.85117055538425e-05 pbeta0 = -7.48385092932104e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.5706062840604e-08 lagidl = -1.97435944398058e-13 wagidl = -8.44806772357702e-15 pagidl = 2.82413559482649e-19
+ bgidl = 2211381960.09463 lbgidl = 698.284479819602 wbgidl = -598.885187811116 pbgidl = -0.00099883030964084
+ cgidl = -2927.80630447562 lcgidl = 0.0131817527583409 wcgidl = 0.00485738171275975 pcgidl = -1.88552582360474e-8
+ egidl = 0.601724962201199 legidl = -6.96926817354889e-06 wegidl = 4.15078228088052e-07 pegidl = 9.96888301105338e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.7070300465303 lkt1 = 2.90346977055966e-07 wkt1 = 1.5881804473722e-07 pkt1 = -4.15314058062717e-13
+ kt2 = -0.019032
+ at = 821473.927825869 lat = -0.995309437347858 wat = -0.686457457785689 pat = 1.423696591039e-6
+ ute = -1.28948672782677 lute = -2.11517772785273e-06 wute = -3.8136522419623e-07 pute = 3.02556291298691e-12
+ ua1 = 2.2096e-11
+ ub1 = -3.77453900358199e-18 lub1 = -9.82679343845922e-24 wub1 = 2.99512763577079e-26 pub1 = 1.40563042951327e-29
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.59 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 1e-06 wmax = 1.5e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.996891024552643+0*(0.0/sqrt(l*w*mult))} lvth0 = -9.54026616871896e-08 wvth0 = 7.47752040531132e-09 pvth0 = 1.157729031243e-13
+ k1 = 0.516366410611791 lk1 = 8.22249534897824e-08 wk1 = 9.30101324024297e-08 pk1 = -1.17615066821505e-13
+ k2 = 0.0572221682158124 lk2 = -6.35548847591476e-08 wk2 = -4.00301076468463e-08 pk2 = 7.9267251225732e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 113831.469866933 lvsat = 0.701700110831397 wvsat = 0.0951485046135199 pvsat = -1.0037160487339e-6
+ ua = 3.37262098104143e-09 lua = 2.48079254106215e-15 wua = -1.00818101788972e-15 pua = -3.43027075265134e-21
+ ub = -1.36597784349008e-18 lub = -8.56055243025542e-25 wub = 1.39377860891751e-24 pub = 1.61320906626607e-30
+ uc = 5.53920772381503e-11 luc = -2.6511659597242e-16 wuc = -9.51749725244217e-17 puc = 3.08881508350703e-22
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0203456249060647 lu0 = 8.45210530891698e-09 wu0 = -1.88135472535131e-09 pu0 = -1.13920617648542e-14
+ a0 = 1.52825156478822 la0 = -1.52851250892156e-06 wa0 = -6.58824905710129e-07 pa0 = 1.64676276217943e-12
+ keta = -0.19822061516783 lketa = 7.43370188809937e-07 wketa = 2.69774450255555e-07 pketa = -1.06332117829487e-12
+ a1 = 0.0
+ a2 = 0.5
+ ags = 1.03869035040999 lags = -3.4995035186676e-06 wags = -1.28888408778119e-06 pags = 5.08612449145869e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0829991830721196+0*(0.009/sqrt(l*w*mult))} lvoff = -7.72211121958313e-08 wvoff = -2.29078346935477e-08 pvoff = 1.1045754221159e-13
+ nfactor = {1.6463159853779+0*(0.02/sqrt(l*w*mult))} lnfactor = -5.58934792695095e-07 wnfactor = 1.61312324770197e-08 pnfactor = 4.1721971208111e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -9.79807366882455e-06 lcit = 2.16107302363897e-11 wcit = 2.11672533643287e-11 pcit = -3.09121181945133e-17
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -0.0639155722424 leta0 = 5.66092622993342e-07 weta0 = 2.05857698028963e-07 peta0 = -8.09742284485414e-13
+ etab = 0.0547604095769366 letab = -4.90745694872928e-07 wetab = -1.78458038421308e-07 petab = 7.01965586420406e-13
+ dsub = 0.0203166040909997 ldsub = 2.12284733622503e-06 wdsub = 7.7196636760861e-07 pdsub = -3.0365335668203e-12
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.48864146385087 lpclm = -7.00477655040517e-06 wpclm = -2.35580605149164e-06 ppclm = 1.00196744063588e-11
+ pdiblc1 = 0.391633981428347 lpdiblc1 = -6.42727411831028e-09 wpdiblc1 = -2.3372568389963e-09 ppdiblc1 = 9.19361146247595e-15
+ pdiblc2 = 0.00129
+ pdiblcb = -0.025
+ drout = 0.700317988756931 ldrout = -5.51941510365332e-07 wdrout = -2.00711693025846e-07 pdrout = 7.89500448075633e-13
+ pscbe1 = 358394901.079153 lpscbe1 = -600.36818684561 wpscbe1 = -200.371488584527 ppscbe1 = 0.00085877025667308
+ pscbe2 = 1.45129969248697e-08 lpscbe2 = 1.694584114615e-15 wpscbe2 = 6.75389186862853e-16 ppscbe2 = -2.42394328505001e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.000632891269690017 lalpha0 = -2.26272379929466e-09 walpha0 = -8.76467569906308e-10 palpha0 = 3.23661369885388e-15
+ alpha1 = -3.65975665303e-10 lalpha1 = 7.07615778741678e-16 walpha1 = 5.23493787503403e-16 palpha1 = -1.01217785560677e-21
+ beta0 = 195.77318687791 lbeta0 = -0.000370391148191962 wbeta0 = -0.00022643889541216 pbeta0 = 5.29809720720671e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -5.1184190781514e-08 lagidl = 6.56772026758113e-14 wagidl = 7.31270969185693e-14 pagidl = -3.84627585130572e-20
+ bgidl = 3159440770.71536 lbgidl = -3030.90959205108 wbgidl = -1689.62555704264 pbgidl = 0.00329160238643321
+ cgidl = -975.11706476352 lcgidl = 0.00550083987048719 wcgidl = 0.00105199815013115 pcgidl = -3.88676296552999e-9
+ egidl = -2.14674585215088 legidl = 3.84185551705908e-06 wegidl = 4.34650737176215e-06 pegidl = -5.4954131827344e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.71996926438635 lkt1 = 3.41243455188831e-07 wkt1 = 1.69029288134732e-07 pkt1 = -4.55480035023045e-13
+ kt2 = -0.019032
+ at = 342067.494632585 lat = 0.890438164650087 wat = 0.0685276089186881 pat = -1.546040943768e-6
+ ute = -2.21996876717829 lute = 1.5448780263467e-06 wute = 7.47291121040287e-07 pute = -1.41401246428265e-12
+ ua1 = -9.30819072264911e-11 lua1 = 4.53052873964938e-16 wua1 = -5.68578961955995e-16 pua1 = 2.23650818974871e-21
+ ub1 = -5.61341139742245e-18 lub1 = -2.59357968292582e-24 wub1 = 3.3507416759954e-24 pub1 = 9.93958654205852e-31
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.60 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 1e-06 wmax = 1.5e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.03977142796045+0*(0.0/sqrt(l*w*mult))} lvth0 = -1.2493187296173e-08 wvth0 = 4.85155487963733e-08 pvth0 = 3.64256700400413e-14
+ k1 = 0.563739228603907 lk1 = -9.37062696206323e-09 wk1 = 2.52477693095996e-08 pk1 = 1.34038010302968e-14
+ k2 = 0.0201881928785313 lk2 = 8.05049172536212e-09 wk2 = 4.72106462594718e-09 pk2 = -7.25936411957574e-15
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 600010.573917718 lvsat = -0.238329617746317 wvsat = -0.560226268304448 pvsat = 2.6345435157686e-7
+ ua = 3.51607403808389e-09 lua = 2.20342533800527e-15 wua = -1.12924954105922e-15 pua = -3.19618415776048e-21
+ ub = -9.15510246684732e-19 lub = -1.72703659378666e-24 wub = 8.46242753185329e-25 pub = 2.67187238100351e-30
+ uc = -1.57967780285461e-10 luc = 1.4741575534877e-16 wuc = 1.26745422581434e-16 puc = -1.20202685188445e-22
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0225037162931251 lu0 = 4.27942482157873e-09 wu0 = -4.17539434377875e-09 pu0 = -6.95652469242666e-15
+ a0 = 0.677561297221496 la0 = 1.16301376870032e-07 wa0 = 2.98507727058817e-07 pa0 = -2.04244669942491e-13
+ keta = 0.233922892293723 lketa = -9.2181443584513e-08 wketa = -3.48366215678495e-07 pketa = 1.31856889991949e-13
+ a1 = 0.0
+ a2 = 0.5
+ ags = -0.778735126888446 lags = 1.44977288163091e-08 wags = 1.33333924196993e-06 pags = 1.60425722682548e-14
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.11162406423013+0*(0.009/sqrt(l*w*mult))} lvoff = -2.18747613524119e-08 wvoff = 1.80373670641578e-08 pvoff = 3.1289789887058e-14
+ nfactor = {1.53513520729782+0*(0.02/sqrt(l*w*mult))} lnfactor = -3.43966202373382e-07 wnfactor = 1.20872975636905e-07 pnfactor = 2.14701027972754e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -2.00141919265091e-06 lcit = 6.53585982343559e-12 wcit = 1.0014872021683e-11 pcit = -9.34893310660121e-18
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.297552470836224 leta0 = -1.32807645639394e-07 weta0 = -3.11188359598961e-07 peta0 = 1.89968853168463e-13
+ etab = -0.199291028424605 letab = 4.64030760243251e-10 wetab = 1.84938662804726e-07 petab = -6.63752383636513e-16
+ dsub = 1.20147320984086 ldsub = -1.60924866775359e-07 wdsub = -9.1756712819563e-07 pdsub = 2.30187894984673e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -2.23826151027487 lpclm = 2.13471398458185e-06 wpclm = 4.40558731516786e-06 ppclm = -3.05351347504413e-12
+ pdiblc1 = 0.274254457644749 lpdiblc1 = 2.20526622014894e-07 wpdiblc1 = 1.65563118258204e-07 ppdiblc1 = -3.15442603289837e-13
+ pdiblc2 = 0.00254538820099779 lpdiblc2 = -2.42729936357023e-09 wpdiblc2 = -1.79571481503644e-09 ppdiblc2 = 3.47202357344704e-15
+ pdiblcb = -0.025
+ drout = 1.04367746391703 ldrout = -1.21582877238475e-06 wdrout = -6.91855146451699e-07 pdrout = 1.73912877099179e-12
+ pscbe1 = 49857795.5715535 lpscbe1 = -3.81015066113741 wpscbe1 = 240.961838356176 ppscbe1 = 5.4500623665949e-6
+ pscbe2 = 1.47822952910737e-08 lpscbe2 = 1.1738943770676e-15 wpscbe2 = 2.90183188054383e-16 ppscbe2 = -1.67914556032377e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -0.000963891669385505 lalpha0 = 8.24663997322561e-10 walpha0 = 1.40758032684495e-09 palpha0 = -1.17960432975418e-15
+ alpha1 = 0.0
+ beta0 = -5.15741572151012 lbeta0 = 1.81091765870305e-05 wbeta0 = 6.09734441296664e-05 pbeta0 = -2.59034748451479e-11
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -6.26003055960495e-08 lagidl = 8.77503177502897e-14 wagidl = 1.28567243720057e-13 pagidl = -1.45656559554467e-19
+ bgidl = 1530396369.85791 lbgidl = 118.855902228801 wbgidl = 124.340428385663 pbgidl = -0.000215709916222345
+ cgidl = 2702.85124598773 lcgidl = -0.00161053024819191 wcgidl = -0.00131646575987761 pcgidl = 6.92673846791489e-10
+ egidl = -2.51709183098972 legidl = 4.55792131887388e-06 wegidl = 4.87625248196911e-06 pegidl = -6.51967800204511e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.55672665497878 lkt1 = 2.56130536862458e-08 wkt1 = -3.42414808281235e-08 pkt1 = -6.24549868795209e-14
+ kt2 = -0.019032
+ at = 1577233.87198086 lat = -1.4977622017847 wat = -1.46323698530671 pat = 1.41563355798979e-6
+ ute = -1.5516114918939 lute = 2.52605892797955e-07 wute = 1.77477476966416e-07 pute = -3.12274934397605e-13
+ ua1 = -2.42589621067018e-10 lua1 = 7.42126786214166e-16 wua1 = 1.13715792391199e-15 pua1 = -1.06154260776146e-21
+ ub1 = -1.00950155823991e-17 lub1 = 6.07162441674749e-24 wub1 = 7.47263443845133e-24 pub1 = -6.97574161146651e-30
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.81e-6
+ sbref = 2.81e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.61 pmos
* DC IV MOS Parameters
+ lmin = 8.0e-07 lmax = 1e-06 wmin = 1e-06 wmax = 1.5e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.33943978089698+0*(0.0/sqrt(l*w*mult))} lvth0 = 2.67248718511838e-07 wvth0 = 4.08575887095996e-07 pvth0 = -2.99692456064349e-13
+ k1 = 0.468398584179135 lk1 = 7.96303413116826e-08 wk1 = 1.84863599598273e-07 pk1 = -1.35598374623331e-13
+ k2 = 0.0177083111486775 lk2 = 1.03654737195893e-08 wk2 = -1.42611334296544e-08 pk2 = 1.04606126763187e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1398883.12328471 lvsat = -0.984081136943155 wvsat = -1.29759835508342 pvsat = 9.51794881445463e-7
+ ua = 2.21337107283139e-08 lua = -1.51762316005079e-14 wua = -2.12517212529349e-14 pua = 1.5588243797634e-20
+ ub = -1.61646720300905e-17 lub = 1.25081321768315e-23 wub = 1.73092211115789e-23 pub = -1.26964002314487e-29
+ uc = 6.69148433481003e-12 luc = -6.29449147057633e-18 wuc = -9.42599740781478e-18 puc = 6.91401622861918e-24
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0685305310464626 lu0 = -3.86868368847355e-08 wu0 = -5.42713809465791e-08 pu0 = 3.98083292812205e-14
+ a0 = 0.824654602913926 la0 = -2.10109594603801e-08 wa0 = 3.72068929027748e-07 pa0 = -2.72914419786498e-13
+ keta = 0.867918192855693 lketa = -6.84019226635616e-07 wketa = -9.66723570875022e-07 pketa = 7.09096572854683e-13
+ a1 = 0.0
+ a2 = 0.5
+ ags = -6.26060756920095 lags = 5.13185306307724e-06 wags = 6.30360710671697e-06 pags = -4.62372733081243e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.323721513545748+0*(0.009/sqrt(l*w*mult))} lvoff = 1.76119268070964e-07 wvoff = 2.40638811141423e-07 pvoff = -1.7650977116629e-13
+ nfactor = {0.131713340025851+0*(0.02/sqrt(l*w*mult))} lnfactor = 9.66135127834338e-07 wnfactor = 1.63768277547341e-06 pnfactor = -1.20124850422363e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -1.3337625e-05 lcit = 1.7118264625625e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.699767444137878 leta0 = -5.08277334291354e-07 weta0 = -5.02635182294822e-07 peta0 = 3.68685419389163e-13
+ etab = -0.91285902253384 letab = 6.66583321101184e-07 wetab = 8.59887070189447e-07 petab = -6.3073146541931e-13
+ dsub = 3.83063293489018 ldsub = -2.61525861590753e-06 wdsub = -3.13182803510794e-06 pdsub = 2.29721152289185e-12
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -4.0010580173615 lpclm = 3.78029333792975e-06 wpclm = 5.29562155800823e-06 ppclm = -3.88436489090683e-12
+ pdiblc1 = 0.717174995843783 lpdiblc1 = -1.92941914996594e-07 wpdiblc1 = -8.04443022901061e-07 ppdiblc1 = 5.90062979513043e-13
+ pdiblc2 = -0.0244746288612415 lpdiblc2 = 2.27960216641154e-08 wpdiblc2 = 8.97857407518224e-09 ppdiblc2 = -6.58582897701655e-15
+ pdiblcb = -0.025
+ drout = -3.21058266826395 ldrout = 2.75554433230685e-06 wdrout = 5.46639266251697e-06 pdrout = -4.00962634991951e-12
+ pscbe1 = -1139361348.97907 lpscbe1 = 1106.33186687259 wpscbe1 = 1151.94571640639 ppscbe1 = -0.000844957942712668
+ pscbe2 = 2.5411980972332e-08 lpscbe2 = -8.74897035481541e-15 wpscbe2 = -7.04129051679537e-15 ppscbe2 = 5.16482180052199e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -0.000494700484325197 lalpha0 = 3.86671680112838e-10 walpha0 = 6.71894716286117e-10 palpha0 = -4.92838133869449e-16
+ alpha1 = 0.0
+ beta0 = -107.541757740489 lbeta0 = 0.000113685471783458 wbeta0 = 0.000155077700585582 pbeta0 = -1.13750268768027e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.18120707494248e-07 lagidl = -8.09536515745681e-14 wagidl = -1.28191973527878e-13 pagidl = 9.40294535425662e-20
+ bgidl = 1177707612.36503 lbgidl = 448.092620792189 wbgidl = -498.187523110941 pbgidl = 0.000365423039139489
+ cgidl = 2692.53677096935 lcgidl = -0.00160090163418987 wcgidl = -0.00268126761191528 pcgidl = 1.96672319967792e-9
+ egidl = 10.4464504590863 legidl = -7.54361022662358e-06 wegidl = -9.83835964432271e-06 pegidl = 7.21648599090893e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.1214205493486 lkt1 = -3.80747372450056e-07 wkt1 = -4.72097902199892e-07 pkt1 = 3.46286171753132e-13
+ kt2 = -0.019032
+ at = -200382.980606 lat = 0.161652018189404 wat = 0.248472580105206 pat = -1.82255879870069e-7
+ ute = -0.551952469712297 lute = -6.8058080270368e-07 wute = -7.32994111310356e-07 pute = 5.37654845616704e-13
+ ua1 = 5.524e-10
+ ub1 = -3.5909e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.41e-6
+ sbref = 2.41e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.62 pmos
* DC IV MOS Parameters
+ lmin = 6e-07 lmax = 8.0e-07 wmin = 1e-06 wmax = 1.5e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.003144025375+0*(0.0/sqrt(l*w*mult))} lvth0 = 2.05741003576901e-8
+ k1 = 0.44254341525 lk1 = 9.85952369970487e-8
+ k2 = 0.060159521830025 lk2 = -2.07727015712325e-8
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 8777.45034400001 lvsat = 0.0355683246872243
+ ua = 1.9726835474425e-09 lua = -3.88017358202812e-16
+ ub = 6.87228769500001e-19 lub = 1.47178680827902e-25
+ uc = 4.14959472645e-13 luc = -1.69062910155397e-18
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.018260895675 lu0 = -1.81380799159088e-9
+ a0 = 0.67330385 la0 = 9.00055745557503e-8
+ keta = -0.0996496058249999 lketa = 2.56965915356666e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.771841104225501 lags = -2.64832011244249e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.093344647362825+0*(0.009/sqrt(l*w*mult))} lvoff = 7.13668484145893e-9
+ nfactor = {1.06762466205+0*(0.02/sqrt(l*w*mult))} lnfactor = 2.79639493573015e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -0.022662087845 leta0 = 2.16283395657467e-08 peta0 = 6.31088724176809e-30
+ etab = -0.0150166811125 letab = 8.01147445692432e-9
+ dsub = 0.247563769959 ldsub = 1.29405319153238e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.293549260715 lpclm = -1.03327573575756e-7
+ pdiblc1 = 0.6023909982125 lpdiblc1 = -1.0874727881406e-7
+ pdiblc2 = 0.00328404983666751 lpdiblc2 = 2.4348920458057e-9
+ pdiblcb = -0.025
+ drout = 0.28951360501675 ldrout = 1.88206215374089e-7
+ pscbe1 = 450011179.51075 lpscbe1 = -59.4808296373326
+ pscbe2 = 1.046761763215e-08 lpscbe2 = 2.21279487702481e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.9926008739325e-05 lalpha0 = -5.4795256824536e-12
+ alpha1 = 0.0
+ beta0 = 45.5070542532001 lbeta0 = 1.42340294202655e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -9.69312851200001e-08 lagidl = 7.67880602679456e-14 wagidl = -1.26217744835362e-29 pagidl = -6.01853107621011e-36
+ bgidl = 2428272495 lbgidl = -469.202973444975
+ cgidl = -706.3914 lcgidl = 0.000892229173857
+ egidl = -2.64167104212725 legidl = 2.0565923351241e-06 pegidl = -2.01948391736579e-28
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.605875525500001 lkt1 = -2.53972251681223e-8
+ kt2 = -0.019032
+ at = 46675.25 lat = -0.01956642925125
+ ute = -1.849518965 lute = 2.71190709422324e-7
+ ua1 = 5.5346701e-10 lua1 = -7.8265717005015e-19
+ ub1 = -8.1825107825e-18 lub1 = 3.36796946701766e-24
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.02e-6
+ sbref = 2.01e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.63 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 6e-07 wmin = 1e-06 wmax = 1.5e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.023/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.945969393690952+0*(0.0/sqrt(l*w*mult))} lvth0 = -9.92885151890959e-09 wvth0 = 1.52125888064328e-07 pvth0 = -8.11599219117587e-14
+ k1 = 0.53554630992352 lk1 = 4.8977727674251e-08 wk1 = 3.5919894534606e-07 pk1 = -1.9163443333685e-13
+ k2 = -0.0147690322045585 lk2 = 1.9202056648988e-08 wk2 = -5.05293798885701e-08 pk2 = 2.69576768174516e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 448557.439887698 lvsat = -0.199056498634287 wvsat = -0.570840163966135 pvsat = 3.04546081676753e-7
+ ua = -4.97704354346501e-09 lua = 3.3196967934318e-15 wua = 5.35678244976655e-15 pua = -2.8578702208627e-21
+ ub = 1.05559583578568e-17 lub = -5.11783789820841e-24 wub = -1.0270147474833e-23 pub = 5.47917502856077e-30
+ uc = -1.7172874972346e-11 luc = 7.69256851402094e-18 wuc = 2.630399338039e-17 puc = -1.4033311988405e-23
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.00474503031703954 lu0 = 5.39697375620783e-09 wu0 = 5.48190899275489e-09 pu0 = -2.92462585717971e-15
+ a0 = 0.193150534030572 la0 = 3.46169769392019e-07 wa0 = 1.09282788672423e-06 pa0 = -5.83029141706812e-13
+ keta = 0.253554419882806 lketa = -1.62739522199577e-07 wketa = -4.57225756787996e-07 pketa = 2.4393222737518e-13
+ a1 = 0.0
+ a2 = 0.5
+ ags = -5.70888775993407 lags = 3.43101805154903e-06 wags = 8.42942134458595e-06 pags = -4.49713843444333e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.202802823126663+0*(0.009/sqrt(l*w*mult))} lvoff = 6.55331689023451e-08 wvoff = 2.48253618259206e-07 pvoff = -1.32444546609378e-13
+ nfactor = {-0.488438775294192+0*(0.02/sqrt(l*w*mult))} lnfactor = 1.10980711771333e-06 wnfactor = 2.93935047023804e-06 pnfactor = -1.56815817262434e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -3.03335653030001e-05 lcit = 2.15181587569771e-11 wcit = 5.76933738108032e-11 pcit = -3.07797033949326e-17
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.621943014343626 leta0 = -3.22271705477396e-07 weta0 = -1.12085532772152e-06 peta0 = 5.97981921616071e-13
+ etab = 0.0848923799799515 letab = -4.5290509181204e-08 wetab = -3.4835259106963e-08 petab = 1.85847849098603e-14
+ dsub = 0.300833217913155 ldsub = -1.54789849154576e-08 wdsub = -5.2728397447393e-08 pdsub = 2.81308636801714e-14
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -1.79901931812534 lpclm = 1.54657322607846e-06 wpclm = 4.54885817394303e-06 ppclm = -2.42683858008948e-12
+ pdiblc1 = 0.878668761349596 lpdiblc1 = -2.56142846836516e-07 wpdiblc1 = 6.25126167119673e-07 ppdiblc1 = -3.33507935789181e-13
+ pdiblc2 = 0.010474118261525 lpdiblc2 = -1.40104540919789e-09 wpdiblc2 = 2.08290722090711e-08 ppdiblc2 = -1.11124141689005e-14
+ pdiblcb = -1.63834261212 lpdiblcb = 8.60726350279083e-07 wpdiblcb = 2.30773495243213e-06 ppdiblcb = -1.2311881357973e-12
+ drout = -0.908418287814499 ldrout = 8.27308869859026e-7
+ pscbe1 = 4029357792.51061 lpscbe1 = -1969.08014440582 wpscbe1 = -5295.28846726259 ppscbe1 = 0.00282506287372693
+ pscbe2 = -5.90866543879953e-08 lpscbe2 = 3.93203467711325e-14 wpscbe2 = 1.04584910706275e-13 ppscbe2 = -5.57965727863514e-20
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -3.51020111327407e-05 lalpha0 = 3.45482980593929e-11 walpha0 = 1.63726078963246e-10 palpha0 = -8.73486817572865e-17
+ alpha1 = 0.0
+ beta0 = -5.75951637511275 lbeta0 = 2.87743747050846e-05 wbeta0 = 9.08616636522264e-05 pbeta0 = -4.8475151866781e-11
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 2.45703134773119e-07 lagidl = -1.06009115917133e-13 wagidl = -4.53204528633383e-14 pagidl = 2.41786882048553e-20
+ bgidl = 3846825916.36753 lbgidl = -1226.00831651166 wbgidl = -4144.6919745681 pbgidl = 0.00221121389189195
+ cgidl = 1372.79068787999 lcgidl = -0.000217024865937417 wcgidl = 0.00230773495243213 pcgidl = -1.2311881357973e-9
+ egidl = -0.400565919934039 legidl = 8.60951546908412e-07 wegidl = 5.84934816729561e-06 pegidl = -3.12065649399304e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.498179608181998 lkt1 = -8.28535355368624e-08 wkt1 = -3.4616024286482e-07 pkt1 = 1.84678220369595e-13
+ kt2 = -0.019032
+ at = -591.602242400084 lat = 0.00565067275433166 wat = 0.0461546990486426 pat = -2.4623762715946e-8
+ ute = -0.885881090824721 lute = -2.4291491463956e-07 wute = -9.09247571258257e-07 pute = 4.85088125504136e-13
+ ua1 = 5.52e-10
+ ub1 = -6.10701479999998e-19 lub1 = -6.71628654912602e-25
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 1.81e-6
+ sbref = 1.81e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.64 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 7.5e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.011588699336+0*(0.0/sqrt(l*w*mult))} wvth0 = 1.65581558424102e-8
+ k1 = 0.62249005992 wk1 = -3.50205375899277e-8
+ k2 = 0.020618136649224 wk2 = 5.37171239304811e-9
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -192534.395056 wvsat = 0.253712779702473
+ ua = 2.0254698305032e-09 wua = 2.1527805622444e-16
+ ub = 8.38826662912e-19 wub = -5.44649124305302e-25
+ uc = -7.9046095641168e-11 wuc = 3.15756663168246e-17
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.01800925453888 wu0 = 1.74418989818813e-10
+ a0 = 1.0051307358728 wa0 = -8.73986513922682e-8
+ keta = -0.0094997103408 wketa = 1.22609864794236e-9
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.20935864688912 wags = -5.78063730952386e-8
+ b0 = 1.32496821192e-07 wb0 = -1.23275837417964e-13
+ b1 = -1.5480597312e-07 wb1 = 1.44032406226687e-13
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.10399611253736+0*(0.009/sqrt(l*w*mult))} wvoff = -3.42763195134506e-9
+ nfactor = {1.5150988704+0*(0.02/sqrt(l*w*mult))} wnfactor = 5.1657192106619e-8
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -8.60812e-06 wcit = 1.266107649672e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -2.39700789405 wpclm = 2.30790850285898e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0092842962121584 wpdiblc2 = -5.43936710852985e-9
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 222315123.63024 wpscbe1 = 2.23528773334283
+ pscbe2 = 1.5010532126536e-08 wpscbe2 = -1.09872821838481e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.000187434197076512 walpha0 = -1.14618162922923e-10
+ alpha1 = 0.0
+ beta0 = 42.721745458408 wbeta0 = -3.42600373690757e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -9.39353920000001e-09 wagidl = 2.73479252329152e-14
+ bgidl = 1026425244.0 wbgidl = 459.597076830936
+ cgidl = 1944.3248 wcgidl = -0.000506443059868801
+ egidl = 2.6925648631184 wegidl = -1.09102167434334e-6
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.52878376 wkt1 = -2.53221529934397e-8
+ kt2 = -0.019032
+ at = -394187.3684 wat = 0.50732933522357
+ ute = -1.9526406168 wute = 3.6894376911442e-7
+ ua1 = 2.2096e-11
+ ub1 = -4.9189672856e-18 wub1 = 1.71405653612595e-24
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.65 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 7.5e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.0233545495998+0*(0.0/sqrt(l*w*mult))} lvth0 = 2.34534635062795e-07 wvth0 = 2.75051735229549e-08 pvth0 = -2.18212431670234e-13
+ k1 = 0.647374860217969 lk1 = -4.96041291163553e-07 wk1 = -5.81735050959592e-08 pk1 = 4.61519793546317e-13
+ k2 = 0.0168011195684362 lk2 = 7.60865290649684e-08 wk2 = 8.92308798711554e-09 pk2 = -7.07913631612211e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -372816.946108396 lvsat = 3.59366313281569 wvsat = 0.421448746896928 pvsat = -3.34356574075052e-6
+ ua = 1.87249812286097e-09 lua = 3.04926229914486e-15 wua = 3.57603850845014e-16 pua = -2.83705193869817e-21
+ ub = 1.22584198659164e-18 lub = -7.71457188964471e-24 wub = -9.04730503548781e-25 pub = 7.17768397355678e-30
+ uc = -1.01483048487816e-10 luc = 4.4724711175342e-16 wuc = 5.24511418670629e-17 puc = -4.16121396258053e-22
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0178853163577864 lu0 = 2.47052235251953e-09 wu0 = 2.89731817137358e-10 pu0 = -2.29858881991832e-15
+ a0 = 1.06723423672922 la0 = -1.23794044483895e-06 wa0 = -1.45180121210086e-07 pa0 = 1.15178721752083e-12
+ keta = -0.010370948251449 lketa = 1.73668252481123e-08 wketa = 2.0367036274377e-09 pketa = -1.61581984117952e-14
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.250434545473801 lags = -8.18786629817225e-07 wags = -9.6023635593817e-08 pags = 7.61803993101726e-13
+ b0 = 2.2009383730957e-07 lb0 = -1.74611555876466e-12 wb0 = -2.04776626795848e-13 pb0 = 1.62459639256799e-18
+ b1 = -2.57152136601449e-07 lb1 = 2.04011776148828e-12 wb1 = 2.39255890806808e-13 pb1 = -1.89813780599526e-18
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.101560514957365+0*(0.009/sqrt(l*w*mult))} lvoff = -4.85499965388215e-08 wvoff = -5.69372655335806e-09 pvoff = 4.51712080796989e-14
+ nfactor = {1.47839244045939+0*(0.02/sqrt(l*w*mult))} lnfactor = 7.31687804753192e-07 wnfactor = 8.58090747619355e-08 pnfactor = -6.80766723669196e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -1.760479400505e-05 lcit = 1.79335246263034e-10 wcit = 2.10316359710626e-11 pcit = -1.66854589134605e-16
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -4.03695536921804 lpclm = 3.26899011959994e-05 wpclm = 3.83372547344017e-06 ppclm = -3.0414880212165e-11
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0131493872004256 lpdiblc2 = -7.70448105400798e-08 wpdiblc2 = -9.03547095455961e-09 ppdiblc2 = 7.16829539953535e-14
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 220726778.827996 lpscbe1 = 31.6612790572453 wpscbe1 = 3.71309326741914 ppscbe1 = -2.94578440025364e-5
+ pscbe2 = 1.50183394402376e-08 lpscbe2 = -1.55627126706972e-16 wpscbe2 = -1.82512536956875e-17 ppscbe2 = 1.44796412451011e-22
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.000268879265917411 lalpha0 = -1.62348568696541e-09 walpha0 = -1.90395143642909e-10 palpha0 = 1.51050082406674e-15
+ alpha1 = 0.0
+ beta0 = 45.1561860661261 lbeta0 = -4.85269340261517e-05 wbeta0 = -5.6910218849721e-06 pbeta0 = 4.51497505795357e-11
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -2.8826355050908e-08 lagidl = 3.87364131928154e-13 wagidl = 4.54283336974951e-14 pagidl = -3.60405912530746e-19
+ bgidl = 699845977.616684 lbgidl = 6509.86943934814 wbgidl = 763.448385749572 pbgidl = -0.00605682158558615
+ cgidl = 2304.191760202 lcgidl = -0.00717340985052137 wcgidl = -0.000841265438842502 pcgidl = 6.67418356538419e-9
+ egidl = 3.46782013774325 legidl = -1.54535548930107e-05 wegidl = -1.81232383338594e-06 pegidl = 1.43780801937866e-11
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.5107904119899 lkt1 = -3.58670492526066e-07 wkt1 = -4.20632719421249e-08 pkt1 = 3.33709178269205e-13
+ kt2 = -0.019032
+ at = -754684.095782354 lat = 7.18596331775979 wat = 0.842737653360477 pat = -6.68586338662361e-6
+ ute = -2.21480369730716 lute = 5.22582907610483e-06 wute = 6.12861872196763e-07 pute = -4.86214272738238e-12
+ ua1 = 2.2096e-11
+ ub1 = -6.13693701240367e-18 lub1 = 2.42784056390896e-23 wub1 = 2.84726287776245e-24 pub1 = -2.25887742770428e-29
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.66 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 7.5e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.02137203099661+0*(0.0/sqrt(l*w*mult))} lvth0 = 2.18806313811767e-07 wvth0 = 1.43904057064272e-08 pvth0 = -1.14166355623962e-13
+ k1 = 0.473725586802238 lk1 = 8.81606087726513e-07 wk1 = 8.48633027297128e-08 pk1 = -6.73263436522691e-13
+ k2 = 0.0565602208575576 lk2 = -2.39342499807782e-07 wk2 = -2.19462601653981e-08 pk2 = 1.74110764753487e-13
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 201652.169987663 lvsat = -0.963890472077979 wvsat = -0.149706037561923 pvsat = 1.18769359752771e-6
+ ua = 3.48874844062584e-09 lua = -9.7732676780943e-15 wua = -8.95074270506333e-16 pua = 7.10107620043335e-21
+ ub = -6.94716659785615e-19 lub = 7.52218973418249e-24 wub = 7.8904444647782e-25 pub = -6.25988806135402e-30
+ uc = -6.73873998406581e-11 luc = 1.76749112732951e-16 wuc = 6.81530510699691e-18 puc = -5.40692571428856e-23
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0214450905472105 lu0 = -2.5770963978147e-08 wu0 = -2.25629808108547e-09 pu0 = 1.7900352107782e-14
+ a0 = 0.927407775028598 la0 = -1.28626511804756e-07 wa0 = 1.20621431462071e-08 pa0 = -9.56950729611473e-14
+ keta = -0.000864598987622624 lketa = -5.8051844168201e-08 wketa = -5.30271136041443e-09 pketa = 4.20690870914047e-14
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.0632636570423841 lags = 6.66134549407861e-07 wags = 7.240445850493e-08 pags = -5.74421133571155e-13
+ b0 = -1.30294227160709e-07 lb0 = 1.03368990265062e-12 wb0 = 1.21226530715687e-13 pb0 = -9.61751287565557e-19
+ b1 = 1.52232517324346e-07 lb1 = -1.20773743735529e-12 wb1 = -1.41638047513676e-13 pb1 = 1.12368615813998e-18
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.150131638791409+0*(0.009/sqrt(l*w*mult))} lvoff = 3.36789257254183e-07 wvoff = 2.97899551100635e-08 pvoff = -2.36338757815464e-13
+ nfactor = {1.38755356317404+0*(0.02/sqrt(l*w*mult))} lnfactor = 1.45235849189091e-06 wnfactor = 1.10909961959549e-07 pnfactor = -8.79904737755885e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 8.31187500000056e-08 lcit = 3.90081019812812e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.515096967587026 lpclm = 4.74921995736775e-06 wpclm = -2.02515589348007e-07 ppclm = 1.60665844067036e-12
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00555042427785825 lpdiblc2 = -1.67584001990768e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 225831961.432888 lpscbe1 = -8.84071266457613 wpscbe1 = -1.34884841028838 ppscbe1 = 1.07010956072661e-5
+ pscbe2 = 1.49553947342761e-08 lpscbe2 = 3.43745012762055e-16 wpscbe2 = 3.23840156103338e-17 ppscbe2 = -2.56918749764662e-22
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.000178211057386117 lalpha0 = -9.04169001241345e-10 walpha0 = -4.72588817080664e-11 palpha0 = 3.74928574325353e-16
+ alpha1 = -3.65975665303e-10 lalpha1 = 2.90346977055968e-15 walpha1 = 2.49012038526153e-16 palpha1 = -1.97553825270743e-21
+ beta0 = 167.314143017482 lbeta0 = -0.00101766769628952 wbeta0 = -8.63735881346982e-05 pbeta0 = 6.8524529333457e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -8.67782128484027e-10 lagidl = 1.65554653855239e-13 wagidl = 6.97233707873229e-15 pagidl = -5.53150710758081e-20
+ bgidl = 2182197338.16069 lbgidl = -5250.37249128451 wbgidl = -571.731640456047 pbgidl = 0.00453583582821625
+ cgidl = 4187.78296034524 lcgidl = -0.0221168900548138 wcgidl = -0.00176300523276516 pcgidl = 1.39868108291686e-8
+ egidl = -1.39012130644165 legidl = 2.30869478441374e-05 wegidl = 2.26830394751097e-06 pegidl = -1.7995600709098e-11
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.5095686709697 lkt1 = -3.68363181018527e-07 wkt1 = -2.49012038526155e-08 pkt1 = 1.97553825270742e-13
+ kt2 = -0.019032
+ at = 436389.897615323 lat = -2.26342816423066 wat = -0.328172965573617 pat = 2.60356186324312e-6
+ ute = -1.699377919625 lute = 1.13669609173453e-6
+ ua1 = 2.2096e-11
+ ub1 = -3.742347383625e-18 lub1 = 5.28091684622586e-24
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.67 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 7.5e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.915490871752255+0*(0.0/sqrt(l*w*mult))} lvth0 = -1.97677755481706e-07 wvth0 = -6.82576701610877e-08 pvth0 = 2.1093026404128e-13
+ k1 = 0.710244310164666 lk1 = -4.87414932132182e-08 wk1 = -8.73750286089623e-08 pk1 = 4.23690098964468e-15
+ k2 = -0.00853083929509638 lk2 = 1.66935107579827e-08 wk2 = 2.11468850593483e-08 pk2 = 4.60366254622076e-15
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -60629.0367152952 lvsat = 0.0677939658941424 wvsat = 0.257467606700664 pvsat = -4.13925968047404e-7
+ ua = 1.3875551181159e-09 lua = -1.50821323803483e-15 wua = 8.38736171371378e-16 pua = 2.81124158255169e-22
+ ub = -6.74763651352524e-19 lub = 7.44370447574588e-24 wub = 7.50668777267574e-25 pub = -6.10893717463718e-30
+ uc = -7.20194494486907e-12 luc = -5.99906750269105e-17 wuc = -3.69371187212074e-17 puc = 1.18031120747475e-22
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.012619342019382 lu0 = 8.94516198480906e-09 wu0 = 5.30722523011567e-09 pu0 = -1.18508046544443e-14
+ a0 = 0.304924421448582 la0 = 2.319914871919e-06 wa0 = 4.79366008415927e-07 pa0 = -1.93383716351891e-12
+ keta = 0.284749802495103 lketa = -1.18151752047251e-06 wketa = -1.79584124160544e-07 pketa = 7.27605895747777e-13
+ a1 = 0.0
+ a2 = 0.5
+ ags = -0.818043760842087 lags = 4.13276168419352e-06 wags = 4.38632469732414e-07 pags = -2.01498084687452e-12
+ b0 = 4.59281381367846e-07 lb0 = -1.28540870137449e-12 wb0 = -4.27318152912932e-13 pb0 = 1.19595196821103e-18
+ b1 = 4.0696804634187e-07 lb1 = -2.20974091442336e-12 wb1 = -3.78645512124754e-13 pb1 = 2.05595620522499e-18
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0161583858099393+0*(0.009/sqrt(l*w*mult))} lvoff = -1.9019520321469e-07 wvoff = -8.50969135110639e-08 pvoff = 2.15569314340083e-13
+ nfactor = {2.44744783111203+0*(0.02/sqrt(l*w*mult))} lnfactor = -2.7167409105145e-06 wnfactor = -7.29246643585094e-07 pnfactor = 2.42485547093698e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 2.09880273376491e-05 lcit = -4.32214604727794e-11 wcit = -7.47631972870047e-12 pcit = 2.94081410344419e-17
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.3152084083636 leta0 = -9.25193450340263e-07 weta0 = -1.46881528270744e-07 peta0 = 5.77759225860611e-13
+ etab = -0.135341242729673 letab = 2.57020104983383e-07 wetab = -1.58632050532402e-09 petab = 6.23979963929459e-15
+ dsub = 0.99725287809022 ldsub = -1.71993638223227e-06 wdsub = -1.36981003337909e-07 pdsub = 5.38815461534682e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -2.40673656985794 lpclm = 1.21899937910984e-05 wpclm = 2.19888304333925e-06 ppclm = -7.83925508799813e-12
+ pdiblc1 = 0.798820210103798 lpdiblc1 = -1.60809634054434e-06 wpdiblc1 = -3.81185767116008e-07 ppdiblc1 = 1.49939612087965e-12
+ pdiblc2 = 0.00323876357863765 lpdiblc2 = -7.66547128038908e-09 wpdiblc2 = -1.81314132614594e-09 ppdiblc2 = 7.13200047210168e-15
+ pdiblcb = -0.025
+ drout = -0.0736252657755578 ldrout = 2.49236815105449e-06 wdrout = 5.19369754650709e-07 pdrout = -2.04294352676733e-12
+ pscbe1 = 56555713.4978228 lpscbe1 = 657.008254969243 wpscbe1 = 80.4615025762682 ppscbe1 = -0.000311100329050109
+ pscbe2 = 1.46403562043997e-08 lpscbe2 = 1.58295064522331e-15 wpscbe2 = 5.56893349032426e-16 ppscbe2 = -2.32007883532714e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -0.00125207486777292 lalpha0 = 4.72186783680135e-09 walpha0 = 8.77316234186034e-10 palpha0 = -3.26189226691967e-15
+ alpha1 = 9.95065011212e-10 lalpha1 = -2.45019053571546e-15 walpha1 = -7.42826624170212e-16 palpha1 = 1.92586408620204e-21
+ beta0 = -370.994859387093 lbeta0 = 0.00109977345621389 wbeta0 = 0.000300885495441077 pbeta0 = -8.38040248206159e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -6.2567109938712e-08 lagidl = 4.08249268293409e-13 wagidl = 8.37178331999413e-14 pagidl = -3.57193863796064e-19
+ bgidl = -1403991040.0986 lbgidl = 8855.9174255403 wbgidl = 2556.21878032953 pbgidl = -0.00776797279169592
+ cgidl = -1450.34097166068 lcgidl = 6.06986223511859e-05 wcgidl = 0.00149414932445171 pcgidl = 1.17477709258324e-9
+ egidl = 5.96054825776877 legidl = -5.82694764003214e-06 wegidl = -3.19656771187175e-06 pegidl = 3.5004992874422e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.678651775160581 lkt1 = 2.96726054731816e-07 wkt1 = 1.3058724825414e-07 pkt1 = -4.14060778533439e-13
+ kt2 = -0.019032
+ at = -242453.663511586 lat = 0.406806377679845 wat = 0.612369601582974 pat = -1.09606702738017e-6
+ ute = -1.53781285957876 lute = 5.0117912021735e-07 wute = 1.12609171674236e-07 pute = -4.42948739826468e-13
+ ua1 = -1.28556633882702e-09 lua1 = 5.14369634808777e-15 wua1 = 5.40915708111725e-16 pua1 = -2.12769464243601e-21
+ ub1 = -4.0906336490374e-18 lub1 = 6.65090261265685e-24 wub1 = 1.93394012223146e-24 pub1 = -7.60716314049805e-30
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.68 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 7.5e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.06762101560684+0*(0.0/sqrt(l*w*mult))} lvth0 = 9.64666383118514e-08 wvth0 = 7.44269722400954e-08 pvth0 = -6.4951205464618e-14
+ k1 = 0.675342539992185 lk1 = 1.87412539241265e-08 wk1 = -7.85886212259233e-08 pk1 = -1.27516616174993e-14
+ k2 = 0.00318405406700051 lk2 = -5.95729413209848e-09 wk2 = 2.05418174010283e-08 pk2 = 5.77356388892079e-15
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -32263.8868233412 lvsat = 0.0129498067523002 wvsat = 0.0280456836157985 pvsat = 2.96624673467997e-8
+ ua = 3.09757248546879e-09 lua = -4.8145403678985e-15 wua = -7.39873185496826e-16 pua = 3.33337324280662e-21
+ ub = 7.98810198120365e-19 lub = 4.5945420699208e-24 wub = -7.48771274584002e-25 pub = -3.20976233718189e-30
+ uc = -7.33026001576778e-11 luc = 6.78152723303313e-17 wuc = 4.79724309994639e-17 puc = -4.61419181851914e-23
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0228976635524932 lu0 = -1.09280240910693e-08 wu0 = -4.5419252375784e-09 pu0 = 7.19257702059457e-15
+ a0 = 1.70345380528592 la0 = -3.84148684377405e-07 wa0 = -6.5598881779937e-07 pa0 = 2.61377069742494e-13
+ keta = -0.410074190889693 lketa = 1.61928144856962e-07 wketa = 2.50812534497855e-07 pketa = -1.0456819575153e-13
+ a1 = 0.0
+ a2 = 0.5
+ ags = 1.25830789049175 lags = 1.18125384581287e-07 wags = -5.6193780365871e-07 pags = -8.0373220421415e-14
+ b0 = -2.65406728692056e-07 lb0 = 1.1577938286688e-13 wb0 = 2.46936012815461e-13 pb0 = -1.07721832495643e-19
+ b1 = -4.4710427195032e-07 lb1 = -5.58387816643825e-13 wb1 = 4.15988497248209e-13 pb1 = 5.19527374932314e-19
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.137153534992131+0*(0.009/sqrt(l*w*mult))} lvoff = 4.37495227048237e-08 wvoff = 4.17901398379482e-08 pvoff = -2.97674377454983e-14
+ nfactor = {0.821846257484736+0*(0.02/sqrt(l*w*mult))} lnfactor = 4.26367860101735e-07 wnfactor = 7.84521294276695e-07 pnfactor = -5.0202240575847e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 5.39471838530182e-06 lcit = -1.30717196468712e-11 wcit = 3.13346124233032e-12 pcit = 8.89407647804904e-18
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -0.361366040256384 leta0 = 3.8296662893872e-07 weta0 = 3.01873376632669e-07 peta0 = -2.89910626544661e-13
+ etab = -0.0129598209221188 letab = 2.03950140113675e-08 wetab = 1.15749893571675e-08 petab = -1.92076587863821e-14
+ dsub = -0.058749622954767 ldsub = 3.21849733550717e-07 wdsub = 2.54951756774421e-07 pdsub = -2.18988489806309e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 6.10601353584104 lpclm = -4.2694511020211e-06 wpclm = -3.35797625338866e-06 ppclm = 2.90496014652177e-12
+ pdiblc1 = 0.195230823722821 lpdiblc1 = -4.4105324402979e-07 wpdiblc1 = 2.3908718140097e-07 ppdiblc1 = 3.00095273557333e-13
+ pdiblc2 = -0.00323655973706599 lpdiblc2 = 4.85459872714047e-09 wpdiblc2 = 3.58384423822572e-09 ppdiblc2 = -3.30309810153874e-15
+ pdiblcb = -0.025
+ drout = -0.0422260160787751 ldrout = 2.43165754476951e-06 wdrout = 3.18475966757276e-07 pdrout = -1.65451438340644e-12
+ pscbe1 = 392416212.253692 lpscbe1 = 7.62030132227483 wpscbe1 = -77.7565678753861 ppscbe1 = -5.18489874148389e-6
+ pscbe2 = 1.66733167601565e-08 lpscbe2 = -2.34778875413521e-15 wpscbe2 = -1.46923453290904e-15 ppscbe2 = 1.59744955504613e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.00204307866503226 lalpha0 = -1.64932799464513e-09 walpha0 = -1.39012291411934e-09 palpha0 = 1.12221266352451e-15
+ alpha1 = -2.721624e-10 walpha1 = 2.532215299344e-16
+ beta0 = 216.534942391516 lbeta0 = -3.6218353174061e-05 wbeta0 = -0.000145290456012842 pbeta0 = 2.46431848097501e-11
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 2.81006771672235e-07 lagidl = -2.56052549670765e-13 wagidl = -1.91126842612819e-13 pagidl = 1.74219691111286e-19
+ bgidl = 3393731289.11871 lbgidl = -420.502686613023 wbgidl = -1609.31756050411 pbgidl = 0.000286112550987621
+ cgidl = -1469.30575282898 lcgidl = 9.73671215639873e-05 wcgidl = 0.00256533414476345 pcgidl = -8.96364113413613e-10
+ egidl = 7.6615498055877 legidl = -9.11584263774777e-06 wegidl = -4.59401676855234e-06 pegidl = 6.20247402577941e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.445280851921239 lkt1 = -1.54497792206062e-07 wkt1 = -1.37931324667677e-07 pkt1 = 1.05121224803759e-13
+ kt2 = -0.019032
+ at = -89984.1429881238 lat = 0.112005797400128 wat = 0.0879526591285213 pat = -8.21042470597704e-8
+ ute = -1.11879418384248 lute = -3.08995584412126e-07 wute = -2.25218343348474e-07 pute = 2.10242449607517e-13
+ ua1 = 2.14237924213404e-09 lua1 = -1.48425357242833e-15 wua1 = -1.08183141622345e-15 pua1 = 1.00989503620167e-21
+ ub1 = 2.09376510357481e-18 lub1 = -5.3066632975126e-24 wub1 = -3.86788024446292e-24 pub1 = 3.61068554760736e-30
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.81e-6
+ sbref = 2.81e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.69 pmos
* DC IV MOS Parameters
+ lmin = 8.0e-07 lmax = 1e-06 wmin = 7.5e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.718109497622233+0*(0.0/sqrt(l*w*mult))} lvth0 = -2.29804111284366e-07 wvth0 = -1.69513536444524e-07 pvth0 = 1.62768479095018e-13
+ k1 = 0.958983830680184 lk1 = -2.46039309139574e-07 wk1 = -2.71579857257782e-07 pk1 = 1.67406622174421e-13
+ k2 = -0.0665737131974406 lk2 = 5.91619303980937e-08 wk2 = 6.41553677141201e-08 pk2 = -3.4939903396102e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -84947.5221662708 lvsat = 0.0621302437631018 wvsat = 0.0829665804280513 pvsat = -2.16064644319225e-8
+ ua = -8.43375492873717e-09 lua = 5.95001142989984e-15 wua = 7.18843219917936e-15 pua = -4.06773947531553e-21
+ ub = 1.18445107880782e-17 lub = -5.71667465930781e-24 wub = -8.75069063754215e-24 pub = 4.26006939773636e-30
+ uc = -5.18840908152206e-12 luc = 4.23033438978454e-18 wuc = 1.62712670610109e-18 puc = -2.87834490081574e-24
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = -0.00541541974626225 lu0 = 1.55023807337355e-08 wu0 = 1.45283753466768e-08 pu0 = -1.06096439263106e-14
+ a0 = 2.54512458986592 la0 = -1.16985257013676e-06 wa0 = -1.22866666965231e-06 pa0 = 7.95974707836475e-13
+ keta = -0.54804428880371 lketa = 2.90723921110186e-07 wketa = 3.50696417835777e-07 pketa = -1.97810300266897e-13
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.73791130323108 lags = 6.03918200772061e-07 wags = -2.07856843307025e-07 pags = -4.10909567314513e-13
+ b0 = -6.59895627003987e-07 lb0 = 4.84036741885559e-13 wb0 = 6.13970850738271e-13 pb0 = -4.50350688870776e-19
+ b1 = -4.87880945015402e-06 lb1 = 3.57863112573523e-12 wb1 = 4.53927358528001e-12 pb1 = -3.32957987117081e-18
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0360947163948571+0*(0.009/sqrt(l*w*mult))} lvoff = -5.05893897498246e-08 wvoff = -2.69708866885486e-08 pvoff = 3.44213243221193e-14
+ nfactor = {2.39475512198098+0*(0.02/sqrt(l*w*mult))} lnfactor = -1.04195042944984e-06 wnfactor = -4.67864876708331e-07 pnfactor = 6.67086346786908e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -7.68538653029999e-05 lcit = 6.37077444690769e-11 wcit = 5.90958910753529e-11 pcit = -4.33471315832267e-17
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.495450021078898 leta0 = -4.16875448398073e-07 weta0 = -3.12537025976208e-07 peta0 = 2.83644556342739e-13
+ etab = 0.0540439871761053 letab = -4.21533758673652e-08 wetab = -3.97252914627451e-08 petab = 2.86814098604105e-14
+ dsub = 0.86895068197294 ldsub = -5.44163139600822e-07 wdsub = -3.76261096900221e-07 pdsub = 3.70251865163237e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 3.10568471931273 lpclm = -1.46862915014784e-06 wpclm = -1.3165345246499e-06 ppclm = 9.99264085535492e-13
+ pdiblc1 = -2.0364100358598 lpdiblc1 = 1.64219465659488e-06 wpdiblc1 = 1.75750901210614e-06 ppdiblc1 = -1.1173590975151e-12
+ pdiblc2 = -0.0606977481554302 lpdiblc2 = 5.84949054216256e-08 wpdiblc2 = 4.26807816052112e-08 ppdiblc2 = -3.98002846183066e-14
+ pdiblcb = -0.025
+ drout = 8.75800860962798 ldrout = -5.78340547950087e-06 wdrout = -5.66925647398135e-06 pdrout = 3.93506378868527e-12
+ pscbe1 = -389474785.164539 lpscbe1 = 737.519456867182 wpscbe1 = 454.246758113964 ppscbe1 = -0.000501812663569172
+ pscbe2 = 2.69071152845847e-08 lpscbe2 = -1.19010908456815e-14 wpscbe2 = -8.43237245172111e-15 ppscbe2 = 8.09757361794679e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.000846489397705791 lalpha0 = -5.3230593064953e-10 walpha0 = -5.75956397094807e-10 palpha0 = 3.62184149049524e-16
+ alpha1 = -2.721624e-10 walpha1 = 2.532215299344e-16
+ beta0 = 211.915943733136 lbeta0 = -3.19064948314699e-05 wbeta0 = -0.000142147661611688 pbeta0 = 2.17093705223012e-11
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -7.21129074245953e-08 lagidl = 7.3586436364522e-14 wagidl = 4.8802523194303e-14 pagidl = -4.9755571516491e-20
+ bgidl = -408955461.283352 lbgidl = 3129.32440832106 wbgidl = 978.053320589959 pbgidl = -0.0021292111033681
+ cgidl = -3409.91853337909 lcgidl = 0.00190893885527142 wcgidl = 0.00299649341798233 pcgidl = -1.29885345075981e-9
+ egidl = -2.9514685878175 legidl = 7.91463097587951e-07 wegidl = 2.62714462443091e-06 pegidl = -5.38516240377427e-13
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.571670075318202 lkt1 = -3.65128202188825e-08 wkt1 = -5.31830417406197e-08 pkt1 = 2.60082789499353e-14
+ kt2 = -0.019032
+ at = -33140.9906059998 lat = 0.0589424304356538 wat = 0.0928696291572658 pat = -8.66942631664535e-8
+ ute = -1.33977425 lute = -1.02709587753753e-7
+ ua1 = 5.524e-10
+ ub1 = -3.5909e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.41e-6
+ sbref = 2.41e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.70 pmos
* DC IV MOS Parameters
+ lmin = 6e-07 lmax = 8.0e-07 wmin = 7.5e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.47813862942981+0*(0.0/sqrt(l*w*mult))} lvth0 = 3.27681057042145e-07 wvth0 = 4.41937829580214e-07 pvth0 = -2.85734155140958e-13
+ k1 = 0.202077215733876 lk1 = 3.09155477456617e-07 wk1 = 2.23731194826998e-07 pk1 = -1.95906511085025e-13
+ k2 = 0.101146177148268 lk2 = -6.38614477699356e-08 wk2 = -3.81342300280256e-08 pk2 = 4.00900279957506e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -265793.52061357 lvsat = 0.194781687854188 wvsat = 0.255462478804748 pvsat = -1.48133068370722e-7
+ ua = -1.09537533828398e-08 lua = 7.79844289597641e-15 wua = 1.20268344785563e-14 pua = -7.61673173924987e-21
+ ub = 2.11823070782528e-17 lub = -1.25659949271323e-23 wub = -1.90687438289335e-23 pub = 1.18284130038879e-29
+ uc = 8.80751116119214e-12 luc = -6.03574308784754e-18 wuc = -7.80848044633439e-18 puc = 4.04272012353145e-24
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0113364205305754 lu0 = 3.21482213147364e-09 wu0 = 6.4425732212235e-09 pu0 = -4.67866763827997e-15
+ a0 = 1.00882048359318 la0 = -4.29658266651764e-08 wa0 = -3.12166688994898e-07 pa0 = 1.23717389524357e-13
+ keta = -0.576393948957584 lketa = 3.11518538581353e-07 wketa = 4.43565797316615e-07 pketa = -2.65930454462989e-13
+ a1 = 0.0
+ a2 = 0.5
+ ags = 5.48093623155175 lags = -2.87511429927579e-06 wags = -4.3813703610351e-06 pags = 2.65038346550662e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.370424404962138+0*(0.009/sqrt(l*w*mult))} lvoff = 1.94643108462719e-07 wvoff = 2.57796668948947e-07 pvoff = -1.74457101575762e-13
+ nfactor = {-3.16597963381468+0*(0.02/sqrt(l*w*mult))} lnfactor = 3.03687631760007e-06 wnfactor = 3.93897083849828e-06 pnfactor = -2.56534968449571e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -2.6300000303e-05 lcit = 2.6626231722252e-11 wcit = 3.3773738081913e-11 pcit = -2.47732057517736e-17
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -0.293175615200877 leta0 = 1.61585398941323e-07 weta0 = 2.51687408933072e-07 peta0 = -1.30216887785393e-13
+ etab = -0.0125592052687803 letab = 6.70039880692063e-09 wetab = -2.28645026985189e-09 petab = 1.21983265121734e-15
+ dsub = -0.123303060605106 ldsub = 1.83659941848887e-07 wdsub = 3.45056724357827e-07 pdsub = -1.58838363318647e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.98042535488794 lpclm = -6.43245780045432e-07 wpclm = -6.39073639275069e-07 ppclm = 5.02343138808626e-13
+ pdiblc1 = 1.13830091435022 lpdiblc1 = -6.86471698938917e-07 wpdiblc1 = -4.98613801434035e-07 ppdiblc1 = 5.37518266830688e-13
+ pdiblc2 = 0.024952719904664 lpdiblc2 = -4.33014115279376e-09 wpdiblc2 = -2.01606606432843e-08 ppdiblc2 = 6.29422747817614e-15
+ pdiblcb = -0.025
+ drout = 4.08053505005326 ldrout = -2.35245523618502e-06 wdrout = -3.52718909859064e-06 pdrout = 2.36384665849931e-12
+ pscbe1 = 1802517950.56324 lpscbe1 = -870.318174752824 wpscbe1 = -1258.38041482786 ppscbe1 = 0.000754407930919523
+ pscbe2 = -7.9273512184306e-10 lpscbe2 = 8.41688792668524e-15 wpscbe2 = 1.04766997644317e-14 ppscbe2 = -5.77232539796235e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.000397370907622689 lalpha0 = -2.02875272581124e-10 walpha0 = -3.32568878590475e-10 palpha0 = 1.83658187289004e-16
+ alpha1 = -9.98162406060001e-10 lalpha1 = 5.32524634445041e-16 walpha1 = 9.28696291572661e-16 palpha1 = -4.95464115035473e-22
+ beta0 = 498.782611675889 lbeta0 = -0.000242324630100819 wbeta0 = -0.000421730298279415 pbeta0 = 2.26784632431262e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -1.51871385064519e-07 lagidl = 1.32089678505794e-13 wagidl = 5.11165986289801e-14 pagidl = -5.14529574182038e-20
+ bgidl = 11408498955.0912 lbgidl = -5538.83749336176 wbgidl = -8355.25657982762 pbgidl = 0.0047168183751377
+ cgidl = -6743.25635283364 lcgidl = 0.00435395881253043 wcgidl = 0.00561673537330614 pcgidl = -3.22081402619959e-9
+ egidl = -11.9906258609176 legidl = 7.42173015319325e-06 wegidl = 8.69832365713146e-06 pegidl = -4.99175641675844e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.173004154045801 lkt1 = -3.28936266801796e-07 wkt1 = -4.02746121229217e-07 pkt1 = 2.82414545570219e-13
+ kt2 = -0.019032
+ at = 146491.490606 lat = -0.0728188926957541 wat = -0.0928696291572661 pat = 4.95464115035473e-8
+ ute = -1.849518965 lute = 2.71190709422326e-7
+ ua1 = 5.53467009999999e-10 lua1 = -7.82657170050939e-19
+ ub1 = -8.1825107825e-18 lub1 = 3.36796946701767e-24
+ uc1 = 4.14042724367564e-10 luc1 = -3.8380115453723e-16 wuc1 = -4.86828170207927e-16 puc1 = 3.57090896988366e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.02e-6
+ sbref = 2.01e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.71 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 6e-07 wmin = 7.5e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.02/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.13879863300177+0*(0.0/sqrt(l*w*mult))} lvth0 = -3.86863527752194e-07 wvth0 = -5.98870630705454e-07 pvth0 = 2.69542362463748e-13
+ k1 = 1.42304661908691 lk1 = -3.42237804079246e-07 wk1 = -4.66536667301417e-07 pk1 = 1.72354844699795e-13
+ k2 = -0.175971150774721 lk2 = 8.39820322636192e-08 wk2 = 9.94540384418212e-08 pk2 = -3.3314001174255e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -637055.783867075 lvsat = 0.392851961611249 wvsat = 0.43922089309465 pvsat = -2.46169101186456e-7
+ ua = 2.05209214046227e-08 lua = -8.99345347650876e-15 wua = -1.83666771257239e-14 pua = 8.59835866919162e-21
+ ub = -3.02011161331531e-17 lub = 1.48473182732688e-23 wub = 2.76504791740496e-23 pub = -1.30965260643186e-29
+ uc = 2.25763122787418e-11 luc = -1.33814673280659e-17 wuc = -1.06788889331456e-17 puc = 5.57409740328765e-24
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0266011653936402 lu0 = -4.9289955766957e-09 wu0 = -1.48531702193247e-08 pu0 = 6.68271796596973e-15
+ a0 = 1.37589174437766 la0 = -2.38800179649998e-07 wa0 = -7.6016318299587e-09 pa0 = -3.87695912984247e-14
+ keta = -0.387036926297392 lketa = 2.10495620207028e-07 wketa = 1.38784275246138e-07 pketa = -1.03327988530779e-13
+ a1 = 0.0
+ a2 = 0.5
+ ags = 10.288763113513 lags = -5.44011397993652e-06 wags = -6.45488901397444e-06 pags = 3.75661603444302e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {0.625000419426156+0*(0.009/sqrt(l*w*mult))} lvoff = -3.36421012472558e-07 wvoff = -5.21939485431392e-07 pvoff = 2.41536035466921e-13
+ nfactor = {9.28942885803053+0*(0.02/sqrt(l*w*mult))} lnfactor = -3.60814638984181e-06 wnfactor = -6.15803624301308e-06 pnfactor = 2.821454078526e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 0.000163267131212 lcit = -7.45087807766581e-11 wcit = -1.22433875830932e-10 pcit = 5.85643373087988e-17
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -1.66739056826605 leta0 = 8.94735947476356e-07 weta0 = 1.00915437354001e-06 peta0 = -5.34329300738019e-13
+ etab = 0.125010442407932 letab = -6.6693696076844e-08 wetab = -7.2161345098331e-08 petab = 3.84984384166851e-14
+ dsub = -0.127874954612656 ldsub = 1.86099070161385e-07 wdsub = 3.46144258519657e-07 pdsub = -1.59418568231654e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 6.05622055034028 lpclm = -2.81770289579523e-06 wpclm = -2.7597041311166e-06 ppclm = 1.63371010935854e-12
+ pdiblc1 = -0.805622157225024 lpdiblc1 = 3.50620979361835e-07 wpdiblc1 = 2.19220054350701e-06 ppdiblc1 = -8.98044640267084e-13
+ pdiblc2 = 0.100012372934268 lpdiblc2 = -4.43748413423526e-08 wpdiblc2 = -6.24778571679769e-08 ppdiblc2 = 2.88706634100823e-14
+ pdiblcb = 3.20168522424 lpdiblcb = -1.72145270055816e-06 wpdiblcb = -2.19545598668424e-06 ppdiblcb = 1.17128674617598e-12
+ drout = -6.08974384306358 ldrout = 3.07343940468728e-06 wdrout = 4.82073638455708e-06 pdrout = -2.08981332638742e-12
+ pscbe1 = -7274048803.85581 lpscbe1 = 3972.07557156351 wpscbe1 = 5221.46885043632 ppscbe1 = -0.00270262405134525
+ pscbe2 = 1.62118639518517e-07 lpscbe2 = -7.84971450008202e-14 wpscbe2 = -1.01225821976108e-13 ppscbe2 = 5.38215284632241e-20
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.000256021714065652 lalpha0 = -1.27464771072477e-10 walpha0 = -1.0713718170369e-10 palpha0 = 6.33892498414203e-17
+ alpha1 = 0.0
+ beta0 = 173.334389527734 lbeta0 = -6.86963763436672e-05 wbeta0 = -7.57683809632176e-05 pbeta0 = 4.2212219733484e-11
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 7.0230695549044e-07 lagidl = -3.23618737071979e-13 wagidl = -4.70147387281658e-13 pagidl = 2.26643985385051e-19
+ bgidl = -6486629779.6248 lbgidl = 4008.3031622529 wbgidl = 5469.61720571734 pbgidl = -0.00265882091381947
+ cgidl = 12634.5864255672 lcgidl = -0.00598421719896031 wcgidl = -0.00817030737268648 pcgidl = 4.1346422140012e-9
+ egidl = 19.0291386450114 legidl = -9.1274693095424e-06 wegidl = -1.2228165538157e-05 pegidl = 6.17263020137394e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -2.127159431514 lkt1 = 7.13615344503874e-07 wkt1 = 1.16945235864221e-06 pkt1 = -5.56361204433588e-13
+ kt2 = -0.019032
+ at = 96208.9544848 lat = -0.0459929082624132 wat = -0.0439091197336848 pat = 2.34257349235195e-8
+ ute = -3.61873838683456 lute = 1.21507811706817e-06 wute = 1.63341925409307e-06 pute = -8.71437339154926e-13
+ ua1 = 5.52e-10
+ ub1 = -6.72697966123008e-18 lub1 = 2.59143633616455e-24 wub1 = 5.69062191748555e-24 pub1 = -3.03597524608813e-30
+ uc1 = -1.15568544873513e-09 luc1 = 4.53656674453921e-16 wuc1 = 9.73656340415854e-16 puc1 = -4.22084891851975e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 1.81e-6
+ sbref = 1.81e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.72 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 7e-07 wmax = 7.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.987253+0*(0.0/sqrt(l*w*mult))}
+ k1 = 0.57102
+ k2 = 0.028513
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 180350.0
+ ua = 2.3418663e-9
+ ub = 3.835e-20
+ uc = -3.2639e-11
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0182656
+ a0 = 0.87668
+ keta = -0.0076977
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.1244
+ b0 = -4.8683e-8
+ b1 = 5.688e-8
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.10903374+0*(0.009/sqrt(l*w*mult))}
+ nfactor = {1.59102+0*(0.02/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.99495
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00129
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 225600350.0
+ pscbe2 = 1.4994384e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.8978653e-5
+ alpha1 = 0.0
+ beta0 = 37.686511
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 3.08e-8
+ bgidl = 1701900000.0
+ cgidl = 1200.0
+ egidl = 1.0890786
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.566
+ kt2 = -0.019032
+ at = 351440.0
+ ute = -1.4104
+ ua1 = 2.2096e-11
+ ub1 = -2.3998e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.73 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 7e-07 wmax = 7.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.982929900900416+0*(0.0/sqrt(l*w*mult))} lvth0 = -8.61745175170271e-8
+ k1 = 0.561876635487499 lk1 = 1.82259302226751e-7
+ k2 = 0.0299154777415204 lk2 = -2.79562970729869e-8
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 246590.7999975 lvsat = -1.32041131795416
+ ua = 2.39807234008572e-09 lua = -1.1203833810787e-15
+ ub = -1.0385014362e-19 lub = 2.83454727384998e-24
+ uc = -2.43950424045908e-11 luc = -1.64330969947877e-16
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0183111383187 lu0 = -9.07738303498019e-10
+ a0 = 0.853861454581374 la0 = 4.54853589194898e-7
+ keta = -0.00737758307324998 lketa = -6.38105235995548e-9
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.109307577760675 lags = 3.00844874169697e-7
+ b0 = -8.08685686595833e-08 lb0 = 6.41571193803648e-13
+ b1 = 9.44848137000001e-08 lb1 = -7.49595741913019e-13
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.109928645975254+0*(0.009/sqrt(l*w*mult))} lvoff = 1.78386127322591e-8
+ nfactor = {1.6045069585+0*(0.02/sqrt(l*w*mult))} lnfactor = -2.6884235469456e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.33056270833333e-05 lcit = -6.58927339937606e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.59751210085156 lpclm = -1.20111746501351e-5
+ pdiblc1 = 0.39
+ pdiblc2 = -0.000130141425952753 lpdiblc2 = 2.83083962149362e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 226183951.850308 lpscbe1 = -11.633230401123
+ pscbe2 = 1.49915153768171e-08 lpscbe2 = 5.71817145597481e-17 wpscbe2 = -2.52435489670724e-29
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -1.0946519926495e-05 lalpha0 = 5.96513584156152e-10 palpha0 = 3.94430452610506e-31
+ alpha1 = 0.0
+ beta0 = 36.7920301283888 lbeta0 = 1.7830138926667e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 3.79401545e-08 lagidl = -1.42328305426522e-13
+ bgidl = 1821894263.125 lbgidl = -2391.90624397353
+ cgidl = 1067.77491666667 lcgidl = 0.00263570935975041
+ egidl = 0.804228350801417 legidl = 5.67806386665123e-6
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.572611254166665 lkt1 = 1.31785467987516e-7
+ kt2 = -0.019032
+ at = 483896.477229166 lat = -2.64032185112998
+ ute = -1.31407402679167 lute = -1.92011426857814e-6
+ ua1 = 2.2096e-11
+ ub1 = -1.95228420545833e-18 lub1 = -8.92055832807532e-24
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.74 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 7e-07 wmax = 7.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.00022229729875+0*(0.0/sqrt(l*w*mult))} lvth0 = 5.10147957711113e-8
+ k1 = 0.598450093537499 lk1 = -1.07896410080229e-7
+ k2 = 0.0243055667754387 lk2 = 1.65499596259775e-8
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -18372.3999924995 lvsat = 0.781675553982501
+ ua = 2.17324817974287e-09 lua = 6.63260219122046e-16
+ ub = 4.6495043086e-19 lub = -1.67803492778996e-24 wub = -7.3468396926393e-40
+ uc = -5.73708727862275e-11 luc = 9.72829452639901e-17
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0181289850439 lu0 = 5.3737561289439e-10
+ a0 = 0.945135636255873 la0 = -2.69270587490653e-7
+ keta = -0.00865805078025 lketa = 3.77754459586728e-9
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.169677266717975 lags = -1.78098355021488e-7
+ b0 = 4.787370597875e-08 lb0 = -3.79806285750942e-13
+ b1 = -5.59344410999999e-08 lb1 = 4.43756168139055e-13
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.106349022074237+0*(0.009/sqrt(l*w*mult))} lvoff = -1.05603513845761e-8
+ nfactor = {1.5505591245+0*(0.02/sqrt(l*w*mult))} lnfactor = 1.59153056083605e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 8.31187500000192e-08 lcit = 3.90081019812813e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.812736302554688 lpclm = 7.11054310953039e-06 wpclm = -2.11758236813575e-22 ppclm = -1.61558713389263e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00555042427785826 lpdiblc2 = -1.67584001990768e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 223849544.449075 lpscbe1 = 6.88680238859524
+ pscbe2 = 1.50029898695488e-08 lpscbe2 = -3.38512308994309e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.000108754171779485 lalpha0 = -3.53132451996697e-10
+ alpha1 = 0.0
+ beta0 = 40.3699536148338 lbeta0 = -1.05553349426628e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 9.37953650000001e-09 lagidl = 8.42575002795677e-14
+ bgidl = 1341917210.62499 lbgidl = 1415.99410192054
+ cgidl = 1596.67525000001 lcgidl = -0.00156032407925125
+ egidl = 1.94362934759575 legidl = -3.36137963842162e-06 wegidl = 3.3881317890172e-21
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.5461662375 lkt1 = -7.80162039625644e-8
+ kt2 = -0.019032
+ at = -45929.4316875008 lat = 1.56305464638994
+ ute = -1.69937791962501 lute = 1.13669609173452e-6
+ ua1 = 2.2096e-11
+ ub1 = -3.742347383625e-18 lub1 = 5.28091684622588e-24
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.75 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 7e-07 wmax = 7.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.0158099020975+0*(0.0/sqrt(l*w*mult))} lvth0 = 1.12328717185025e-7
+ k1 = 0.58182829295 lk1 = -4.25144743602903e-8
+ k2 = 0.0225489646151401 lk2 = 2.34595630065237e-8
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 317773.867875 lvsat = -0.540557471405652
+ ua = 2.62025467010599e-09 lua = -1.09504204575379e-15
+ ub = 4.28502306425e-19 lub = -1.53466604808427e-24 wub = 2.75506488473974e-40 pub = 5.25486924121806e-46
+ uc = -6.14888247213663e-11 luc = 1.13480929790618e-16
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.02041942789475 lu0 = -8.47209279313856e-9
+ a0 = 1.00945378835 la0 = -5.22266360343666e-7
+ keta = 0.02081308800325 lketa = -1.12147327164724e-07 pketa = -5.04870979341448e-29
+ a1 = 0.0
+ a2 = 0.5
+ ags = -0.173380912877175 lags = 1.17132270970693e-06 pags = 8.07793566946316e-28
+ b0 = -1.687526937475e-07 lb0 = 4.7229474070426e-13 pb0 = 3.85185988877447e-34
+ b1 = -1.49531326275e-07 lb1 = 8.11919983959343e-13 pb1 = -7.70371977754894e-34
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.141226232817555+0*(0.009/sqrt(l*w*mult))} lvoff = 1.26629331460316e-07 wvoff = 2.11758236813575e-22
+ nfactor = {1.3756662131+0*(0.02/sqrt(l*w*mult))} lnfactor = 8.47095197540078e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.0993350499999996 leta0 = -7.60545158502511e-8
+ etab = -0.137672675 letab = 2.66190805475875e-7
+ dsub = 0.795930427468225 ldsub = -9.28033516098403e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.824985436325498 lpclm = 6.68556461036471e-7
+ pdiblc1 = 0.23858739746545 lpdiblc1 = 5.95582229132667e-7
+ pdiblc2 = 0.000573970313813503 lpdiblc2 = 2.81650635076303e-9
+ pdiblcb = -0.025
+ drout = 0.689698036268675 ldrout = -5.10167874153015e-7
+ pscbe1 = 174810847.309499 lpscbe1 = 199.780762780594
+ pscbe2 = 1.54588283357925e-08 lpscbe2 = -1.82689411706142e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.73262165591325e-05 lalpha0 = -7.21702329976654e-11
+ alpha1 = -9.66752500000001e-11 lalpha1 = 3.80272579251249e-16
+ beta0 = 71.2197822255274 lbeta0 = -0.000131903290031969
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 6.0473887936e-08 lagidl = -1.16722386565696e-13
+ bgidl = 2352911133.5 lbgidl = -2560.75554867792 wbgidl = 3.63797880709171e-12
+ cgidl = 745.626324999994 lcgidl = 0.00178728112248088
+ egidl = 1.26251838755635 legidl = -6.8222627155184e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.486726294999997 lkt1 = -3.11823514986026e-7
+ kt2 = -0.019032
+ at = 657552.511600001 lat = -1.20409509494116
+ ute = -1.37230995149999 lute = -1.49827396224981e-7
+ ua1 = -4.9057671776e-10 lua1 = 2.01660069867255e-15 wua1 = -3.45126646034193e-31 pua1 = 9.4039548065783e-37
+ ub1 = -1.24830109725e-18 lub1 = -4.52942669146163e-24
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.76 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 7e-07 wmax = 7.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.95823489579+0*(0.0/sqrt(l*w*mult))} lvth0 = 1.00715461444446e-9
+ k1 = 0.55984
+ k2 = 0.0333745835465 lk2 = 2.52817467464459e-9
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 8955.15535999998 lvsat = 0.0565450533356633
+ ua = 2.01017292477e-09 lua = 8.45540592620761e-17
+ ub = -3.01666979599998e-19 lub = -1.22880082708501e-25
+ uc = -2.7970035e-12
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.016222347289 lu0 = -3.57016456517949e-10
+ a0 = 0.73934
+ keta = -0.0414523173349999 lketa = 8.24314538380926e-9
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.43242187
+ b0 = 9.75177793449998e-08 lb0 = -4.25405503724543e-14
+ b1 = 1.6427848665e-07 lb1 = 2.05167141619792e-13
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.075734118+0*(0.009/sqrt(l*w*mult))}
+ nfactor = {1.9748656228+0*(0.02/sqrt(l*w*mult))} lnfactor = -3.11459857111921e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.082300500945 leta0 = -4.31181300796619e-8
+ etab = 0.0040520651535 letab = -7.83468823461803e-9
+ dsub = 0.31595571
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.1707598
+ pdiblc1 = 0.54661982
+ pdiblc2 = 0.0020306546
+ pdiblcb = -0.025
+ drout = 0.42584153
+ pscbe1 = 278136550.0
+ pscbe2 = 1.4513967e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 3.0
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.056e-10
+ bgidl = 1028500000.0
+ cgidl = 2300.9933697 lcgidl = -0.00122002883528179
+ egidl = 0.90967406
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.648
+ kt2 = -0.019032
+ at = 39280.8239999999 lat = -0.00866369560811997
+ ute = -1.4498
+ ua1 = 5.524e-10
+ ub1 = -3.5909e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.81e-6
+ sbref = 2.81e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.77 pmos
* DC IV MOS Parameters
+ lmin = 8.0e-07 lmax = 1e-06 wmin = 7e-07 wmax = 7.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.967245361274998+0*(0.0/sqrt(l*w*mult))} lvth0 = 9.41846919701758e-9
+ k1 = 0.55984
+ k2 = 0.0277161192175002 lk2 = 7.81037941808764e-9
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 36989.3514475003 lvsat = 0.0303749911170015
+ ua = 2.13116101730002e-09 lua = -2.83889300551436e-17
+ ub = -1.01647315025e-18 lub = 5.44395051624126e-25
+ uc = -2.7970035e-12
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0159370894125 lu0 = -9.07268025158959e-11
+ a0 = 0.73934
+ keta = -0.032622
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.43242187
+ b0 = 2.42463921175e-07 lb0 = -1.77848498501469e-13
+ b1 = 1.7926096515e-06 lb1 = -1.31488814242351e-12
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.075734118+0*(0.009/sqrt(l*w*mult))}
+ nfactor = {1.707129091775+0*(0.02/sqrt(l*w*mult))} lnfactor = -6.15264667174278e-8
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.036111
+ etab = -0.0043407
+ dsub = 0.31595571
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.1707598
+ pdiblc1 = 0.54661982
+ pdiblc2 = 0.0020306546
+ pdiblcb = -0.025
+ drout = 0.42584153
+ pscbe1 = 278136550.0
+ pscbe2 = 1.4513967e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 3.0
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -3.8731536e-10 lagidl = 4.601389531368e-16 pagidl = -3.76158192263132e-37
+ bgidl = 1028500000.0
+ cgidl = 994.06
+ egidl = 0.90967406
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.649833762500002 lkt1 = 1.71182646256283e-9
+ kt2 = -0.019032
+ at = 103350.5 lat = -0.0684730585025
+ ute = -1.33977425 lute = -1.02709587753742e-7
+ ua1 = 5.524e-10
+ ub1 = -3.5909e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.41e-6
+ sbref = 2.41e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.78 pmos
* DC IV MOS Parameters
+ lmin = 6e-07 lmax = 8.0e-07 wmin = 7e-07 wmax = 7.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.014/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.828617858624995+0*(0.0/sqrt(l*w*mult))} lvth0 = -9.22654971342687e-8
+ k1 = 0.530897353749999 lk1 = 2.12295757376049e-8
+ k2 = 0.0450998900372996 lk2 = -4.94070339708957e-9
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 109662.425989999 lvsat = -0.0229310724252949
+ ua = 6.72221431667525e-09 lua = -3.39594948041338e-15
+ ub = -6.84323036400001e-18 lub = 4.81835060169581e-24 pub = -2.10194769648723e-45
+ uc = -2.66869634775751e-12 luc = -9.41139377056229e-20
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0208051395325 lu0 = -3.66146590578642e-9
+ a0 = 0.550025750749988 la0 = 1.38862948396119e-7
+ keta = 0.0755194635000005 lketa = -7.93223041845675e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = -0.958410806885759 lags = 1.02018272265908e-06 pags = -8.07793566946316e-28
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {0.00846212594580109+0*(0.009/sqrt(l*w*mult))} lvoff = -6.17583659154639e-8
+ nfactor = {2.62316807872499+0*(0.02/sqrt(l*w*mult))} lnfactor = -7.33445643840184e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 2.3337625e-05 lcit = -9.78321462562497e-12
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.0767320706999999 leta0 = -2.97957584638035e-8
+ etab = -0.0159196257675 letab = 8.49319994509009e-9
+ dsub = 0.383830510171498 ldsub = -4.97865052997976e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.04117196900499 lpclm = 9.50533219739843e-8
+ pdiblc1 = 0.405482859491748 lpdiblc1 = 1.03524666217604e-7
+ pdiblc2 = -0.00467761939758253 lpdiblc2 = 4.92055251859675e-9
+ pdiblcb = -0.025
+ drout = -1.1034126202945 ldrout = 1.12171556551177e-06 pdrout = -8.07793566946316e-28
+ pscbe1 = -46937249.4612522 lpscbe1 = 238.443257273825
+ pscbe2 = 1.4604982953e-08 lpscbe2 = -6.67606566052533e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -9.14091422159001e-05 lalpha0 = 6.70491362115737e-11 walpha0 = -2.55125505357527e-26 palpha0 = -2.32937841349906e-32
+ alpha1 = 3.667525e-10 lalpha1 = -1.956642925125e-16
+ beta0 = -121.038933518325 lbeta0 = 9.09831779303589e-05 wbeta0 = -5.42101086242752e-20 pbeta0 = -3.87740912134232e-26
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -7.67447715000002e-08 lagidl = 5.64687148191075e-14 wagidl = -3.94430452610506e-29 pagidl = 2.33218079203142e-35
+ bgidl = -871311305.000008 lbgidl = 1393.52109127403
+ cgidl = 1511.71990149999 lcgidl = -0.000379706126049758
+ egidl = 0.793393764322992 legidl = 8.52921782805594e-8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.764924450499993 lkt1 = 8.61314215640022e-8
+ kt2 = -0.019032
+ at = 10000.0
+ ute = -1.84951896499999 lute = 2.71190709422326e-7
+ ua1 = 5.53467009999997e-10 lua1 = -7.82657170050939e-19
+ ub1 = -8.18251078249996e-18 lub1 = 3.36796946701766e-24
+ uc1 = -3.014538618e-10 luc1 = 1.41019168899609e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.02e-6
+ sbref = 2.01e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.79 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 6e-07 wmin = 7e-07 wmax = 7.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.01896522574999+0*(0.0/sqrt(l*w*mult))} lvth0 = 9.28577496375104e-9
+ k1 = 0.737372672499994 lk1 = -8.8926039192109e-8
+ k2 = -0.0298024831824004 lk2 = 3.50200872274864e-8
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 8471.87622799911 lvsat = 0.0310545918254808
+ ua = -6.47278106967052e-09 lua = 3.64364653317902e-15 wua = -3.15544362088405e-30 pua = -1.50463276905253e-36
+ ub = 1.0437089841e-17 lub = -4.40078662927271e-24
+ uc = 6.88143461284007e-12 luc = -5.18915655583921e-18
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.00477130172499995 lu0 = 4.89266673370393e-9
+ a0 = 1.36471954449999 la0 = -2.95780264038476e-7
+ keta = -0.1830641876 lketa = 5.86333665955381e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.801943458814989 lags = 8.10249201364074e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1420996435236+0*(0.009/sqrt(l*w*mult))} lvoff = 1.85670909053079e-8
+ nfactor = {0.238896906499988+0*(0.02/sqrt(l*w*mult))} lnfactor = 5.38574947897716e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -1.66752500000001e-05 lcit = 1.156385425125e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -0.184225555700001 leta0 = 1.09426440008728e-7
+ etab = 0.018954139115 letab = -1.01121279885481e-8
+ dsub = 0.380856976792497 ldsub = -4.8200110374433e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.00025377297999 lpclm = -4.1662161585569e-7
+ pdiblc1 = 2.4162785072415 lpdiblc1 = -9.69244865835125e-7
+ pdiblc2 = 0.00818799577125495 lpdiblc2 = -1.94331750205389e-9
+ pdiblcb = -0.025
+ drout = 0.995344155215491 ldrout = 2.01833199330351e-9
+ pscbe1 = 400000000.0
+ pscbe2 = 1.33459626518999e-08 lpscbe2 = 6.04932969132978e-16
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 9.85610483694496e-05 lalpha0 = -3.43009103166634e-11
+ alpha1 = 0.0
+ beta0 = 61.9767869151497 lbeta0 = -6.65662399950231e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.1326295e-08 lagidl = 9.48236048602486e-15
+ bgidl = 1552125324.99998 lbgidl = 100.605531985871
+ cgidl = 626.597999999991 lcgidl = 9.25108340100005e-5
+ egidl = 1.05727252660999 legidl = -5.54884607933673e-8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.408402749999993 lkt1 = -1.0407468826125e-7
+ kt2 = -0.019032
+ at = 31675.25 lat = -0.01156385425125
+ ute = -1.21808457999998 lute = -6.56826921471037e-8
+ ua1 = 5.52e-10
+ ub1 = 1.63658843999998e-18 lub1 = -1.8705690636822e-24
+ uc1 = 2.75307723600001e-10 luc1 = -1.66686020719218e-16 wuc1 = -1.97215226305253e-31 puc1 = 9.4039548065783e-38
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 1.81e-6
+ sbref = 1.81e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.80 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 4.2e-07 wmax = 7.0e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.96208759195+0*(0.0/sqrt(l*w*mult))} wvth0 = -1.58644242271684e-8
+ k1 = 0.5312364045 wk1 = 2.5079817304773e-8
+ k2 = 0.0343945296694 wk2 = -3.70775159276777e-9
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 372611.51495 wvsat = -0.12120281259357
+ ua = 3.28797676653e-09 wua = -5.96433714763311e-16
+ ub = -7.252973045e-19 wub = 4.81407842640627e-25
+ uc = -2.128494080165e-11 wuc = -7.15766704299503e-18
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.020397194785 wu0 = -1.34377014203271e-9
+ a0 = 0.8420523785 wa0 = 2.18294603593289e-8
+ keta = -0.0120702663 wketa = 2.7564920309178e-9
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.1451569126205 wags = -1.30852822574389e-8
+ b0 = -6.545243e-08 wb0 = 1.057154928858e-14
+ b1 = 8.045856945e-08 wb1 = -1.48640716526967e-14
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.092582553735+0*(0.009/sqrt(l*w*mult))} wvoff = -1.03709265285736e-8
+ nfactor = {1.161422244+0*(0.02/sqrt(l*w*mult))} wnfactor = 2.70821002968936e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 2.23995210552104e-05 wcit = -7.816732470331e-12
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.1355449946875 wpclm = -7.19037928220968e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00129
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 226351658.0075 wpscbe1 = -0.473629075776046
+ pscbe2 = 1.49873558568e-08 wpscbe2 = 4.43058364213989e-18
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 4.272936315185e-05 walpha0 = -1.49725901839872e-11
+ alpha1 = -1.25145e-10 walpha1 = 7.889215887e-17
+ beta0 = 81.09494519095 wbeta0 = -2.736493736458e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 5.683016e-08 wagidl = -1.640956904496e-14
+ bgidl = 2272060620.0 wbgidl = -359.43267581172
+ cgidl = 949.71 wcgidl = 0.00015778431774
+ egidl = -0.0508939860300006 wegidl = 7.18645558068828e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.5788523915 wkt1 = 8.10222471594909e-9
+ kt2 = -0.019032
+ at = 732681.728 wat = -0.240337072781568
+ ute = -1.36735012 wute = -2.713890265128e-8
+ ua1 = -8.344764728e-10 wua1 = 5.39988426287957e-16
+ ub1 = -1.46721946e-18 wub1 = -5.87904367899239e-25
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.81 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 4.2e-07 wmax = 7.0e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.95671870298142+0*(0.0/sqrt(l*w*mult))} lvth0 = -1.07020775099642e-07 wvth0 = -1.65236964353232e-08 pvth0 = 1.31416058576159e-14
+ k1 = 0.471367267148729 lk1 = 1.19340174873724e-06 wk1 = 5.7057648856971e-08 pk1 = -6.37430265134897e-13
+ k2 = 0.0473883313407055 lk2 = -2.59012010583976e-07 wk2 = -1.10149917460479e-08 pk2 = 1.45658908131609e-13
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 565961.289127783 lvsat = -3.85413869032171 wvsat = -0.201333072570665 pvsat = 1.59727693790474e-6
+ ua = 3.93667753899217e-09 lua = -1.29308800913785e-14 wua = -9.69945949021825e-16 pua = 7.44540798915326e-21
+ ub = -1.43410375157329e-18 lub = 1.41289968567676e-23 wub = 8.38599855975399e-25 pub = -7.12008878376875e-30
+ uc = 5.68668503003855e-12 luc = -5.37639038374093e-16 wuc = -1.8963701465155e-17 puc = 2.35335646184297e-22
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0222445529303648 lu0 = -3.68243228274196e-08 wu0 = -2.47964817168115e-09 pu0 = 2.26420303833873e-14
+ a0 = 0.770531216861796 la0 = 1.42566743312094e-06 wa0 = 5.25318818398487e-08 pa0 = -6.12006872094049e-13
+ keta = -0.0121347915489594 lketa = 1.2862143727588e-09 wketa = 2.99897276633807e-09 pketa = -4.83349095190365e-15
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.120523238094496 lags = 4.91035474332463e-07 wags = -7.07041956840308e-09 pags = -1.19897295486209e-13
+ b0 = -1.24428090398605e-07 lb0 = 1.17559162143389e-12 wb0 = 2.74601838614094e-14 pb0 = -3.36649681700668e-19
+ b1 = 2.47075297756464e-07 lb1 = -3.32125538678055e-12 wb1 = -9.61939566920996e-14 pb1 = 1.62118967008236e-18
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0987156755477492+0*(0.009/sqrt(l*w*mult))} lvoff = 1.22254614320047e-07 wvoff = -7.06872383532163e-09 pvoff = -6.5824473896951e-14
+ nfactor = {1.06461312066773+0*(0.02/sqrt(l*w*mult))} lnfactor = 1.92974514398942e-06 wnfactor = 3.40352314732491e-07 pnfactor = -1.38600275069537e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 3.18343731559181e-05 lcit = -1.88069671523717e-10 wcit = -1.16806326966339e-11 pcit = 7.70210744805101e-17
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 3.4921832298084 lpclm = -2.70425550429736e-05 wpclm = -1.19441204772116e-06 ppclm = 9.47587238792775e-12
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00169355319733023 lpdiblc2 = -8.04422967674809e-09 wpdiblc2 = -1.14966803268533e-09 ppdiblc2 = 2.29169134778732e-14
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 227665608.393377 lpscbe1 = -26.1916365866255 wpscbe1 = -0.934045174689572 ppscbe1 = 9.17770660977283e-6
+ pscbe2 = 1.49808972951348e-08 lpscbe2 = 1.28741771245642e-16 wpscbe2 = 6.69370240098675e-18 ppscbe2 = -4.51118890951127e-23
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -2.46456674335072e-05 lalpha0 = 1.34302050904837e-09 walpha0 = 8.6360247833055e-12 palpha0 = -4.70602444493603e-16
+ alpha1 = -1.25145e-10 walpha1 = 7.889215887e-17
+ beta0 = 79.0810662325608 lbeta0 = 4.01436662864449e-05 wbeta0 = -2.66592620942867e-05 pbeta0 = -1.4066581528768e-11
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.22547785010275e-07 lagidl = -1.30998260673044e-12 wagidl = -5.33371579194604e-14 pagidl = 7.36096277467798e-19
+ bgidl = 2586651225.8371 lbgidl = -6270.89341440686 wbgidl = -482.107377835484 pbgidl = 0.00244533678616421
+ cgidl = 722.337895357603 lcgidl = 0.00453232298474972 wcgidl = 0.000217765570855361 pcgidl = -1.19563660888131e-9
+ egidl = -0.692220079588151 legidl = 1.27838768925719e-05 wegidl = 9.43370069208165e-07 pegidl = -4.47954716641853e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.585687034325392 lkt1 = 1.36238386933169e-07 wkt1 = 8.24305026674155e-09 pkt1 = -2.80714682085171e-15
+ kt2 = -0.019032
+ at = 1117186.80150389 lat = -7.66453380521509 wat = -0.399230020164729 pat = 3.16729336112698e-6
+ ute = -1.24256277693922 lute = -2.48744912683883e-06 wute = -4.50811209744836e-08 pute = 3.57651298656669e-13
+ ua1 = -1.4007783057851e-09 lua1 = 1.12883804193176e-14 wua1 = 8.9698849961276e-16 pua1 = -7.11626274662033e-21
+ ub1 = -4.03150967375607e-19 lub1 = -2.12106146180708e-23 wub1 = -9.76582888086778e-25 pub1 = 7.74772522555089e-30
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.82 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 4.2e-07 wmax = 7.0e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.991554154090468+0*(0.0/sqrt(l*w*mult))} lvth0 = 1.69346450451242e-07 wvth0 = -5.46444948736062e-09 pvth0 = -7.45969851002804e-14
+ k1 = 0.695657642346321 lk1 = -5.86007064344727e-07 wk1 = -6.12802220143735e-08 pk1 = 3.01403825112268e-13
+ k2 = -0.00673640938739918 lk2 = 1.70386890606146e-07 wk2 = 1.956904802491e-08 pk2 = -9.69797243114839e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -92358.8500212175 lvsat = 1.36864742521758 wvsat = 0.0466415020168037 pvsat = -3.70030589457822e-7
+ ua = 1.99743254643039e-09 lua = 2.45412975333539e-15 wua = 1.10835230133993e-16 pua = -1.12897489958532e-21
+ ub = 1.18985521774477e-18 lub = -6.68819474611204e-24 wub = -4.56984327080879e-25 pub = 3.15843481042915e-30
+ uc = -8.46567301618824e-11 luc = 1.79100897768088e-16 wuc = 1.72011682047571e-17 puc = -5.15785281662987e-23
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0179490879805956 lu0 = -2.74623017110095e-09 wu0 = 1.13408188089486e-10 pu0 = 2.07000478786518e-15
+ a0 = 0.940504393683915 la0 = 7.71843849367854e-08 wa0 = 2.91956310481919e-09 pa0 = -2.18407293348098e-13
+ keta = -0.012930246771844 lketa = 7.59696236079017e-09 wketa = 2.69321798627684e-09 pketa = -2.40778387551398e-15
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.227703471939391 lags = -3.59279446777178e-07 wags = -3.65800679288121e-08 pags = 1.14217647329337e-13
+ b0 = 1.40920223016125e-07 lb0 = -9.2955054978344e-13 wb0 = -5.86570826194636e-14 pb0 = 3.4656208251167e-19
+ b1 = -3.96046256902448e-07 lb1 = 1.7809526827137e-12 wb1 = 2.14408529352758e-13 pb1 = -8.42976705966946e-19
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.105413395570451+0*(0.009/sqrt(l*w*mult))} lvoff = 1.7539100960875e-07 wvoff = -5.89824561746087e-10 pvoff = -1.17224853678359e-13
+ nfactor = {0.676394825372468+0*(0.02/sqrt(l*w*mult))} lnfactor = 5.00967693080586e-06 wnfactor = 5.51078419155791e-07 pnfactor = -3.05779935376814e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.3512822984375e-07 lcit = 6.34164465935185e-11 wcit = -3.27870881503779e-14 pcit = -1.5387166893622e-17
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.442100486773002 lpclm = 4.17010449394351e-06 wpclm = -2.33651042083669e-07 ppclm = 1.85367014589766e-12
+ pdiblc1 = 0.39
+ pdiblc2 = 7.9340408009311e-05 lpdiblc2 = 4.76213555839335e-09 wpdiblc2 = 3.44900409805599e-09 ppdiblc2 = -1.35666748647237e-14
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 222411578.98041 lpscbe1 = 15.4912320312974 wpscbe1 = 0.906502059239529 ppscbe1 = -5.42428407333969e-6
+ pscbe2 = 1.50067450789038e-08 lpscbe2 = -7.63217505246486e-17 wpscbe2 = -2.36730650869231e-18 ppscbe2 = 2.67736703948978e-23
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.000272002842532257 lalpha0 = -1.01044192800757e-09 walpha0 = -1.02912941534572e-10 palpha0 = 4.14371837534107e-16
+ alpha1 = -2.4820962080625e-10 lalpha1 = 9.76333784489489e-16 walpha1 = 1.56472834213985e-16 palpha1 = -6.15486675744881e-22
+ beta0 = 128.933774847316 lbeta0 = -0.000355363046772258 wbeta0 = -5.58311642878841e-05 pbeta0 = 2.17368850383648e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -7.42370136578688e-08 lagidl = 2.5121057742727e-13 wagidl = 5.27123749188214e-14 pagidl = -1.05248221552375e-19
+ bgidl = 1746386822.31116 lbgidl = 395.348432288178 wbgidl = -254.980070024627 pbgidl = 0.000643421154010239
+ cgidl = 1385.69707231469 lcgidl = -0.000730440362435185 wcgidl = 0.000133001909081887 pcgidl = -5.23163674383148e-10
+ egidl = 1.04752362259422 legidl = -1.01838846741051e-06 wegidl = 5.64910425675312e-07 pegidl = -1.47703569215243e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.570987199580625 lkt1 = 1.96171744863871e-08 wkt1 = 1.56472834213986e-08 pkt1 = -6.1548667574488e-14
+ kt2 = -0.019032
+ at = -208116.295448057 lat = 2.84976494096864 wat = 0.102243572035838 pat = -8.11149889964179e-7
+ ute = -1.738758598283 lute = 1.44912290277117e-06 wute = 2.48258161100751e-08 pute = -1.96955736238361e-13
+ ua1 = 2.2096e-11
+ ub1 = -3.742347383625e-18 lub1 = 5.28091684622586e-24
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.83 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 4.2e-07 wmax = 7.0e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.012/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.01655284867949+0*(0.0/sqrt(l*w*mult))} lvth0 = 2.67678940610617e-07 wvth0 = 4.68357982962385e-10 pvth0 = -9.79337129488326e-14
+ k1 = 0.572126683685112 lk1 = -1.0009742079607e-07 wk1 = 6.11595269024089e-09 pk1 = 3.63006349307947e-14
+ k2 = 0.0194649940911585 lk2 = 6.73235390162218e-08 wk2 = 1.94415352214109e-09 pk2 = -2.76521136603697e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 577838.667786416 lvsat = -1.26757786206634 wvsat = -0.163946410252956 pvsat = 4.5831801639484e-7
+ ua = 3.05751758831093e-09 lua = -1.71572005932694e-15 wua = -2.75653167213896e-16 pua = 3.91279143824588e-22
+ ub = 1.70795260731809e-19 lub = -2.67971730990178e-24 wub = 1.62460067847262e-25 pub = 7.2184718575733e-31
+ uc = -8.47701696314647e-11 luc = 1.79547112488887e-16 wuc = 1.46766995193955e-17 puc = -4.16485179700854e-23
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0210256991038743 lu0 = -1.48480954075733e-08 wu0 = -3.82197007859201e-10 pu0 = 4.01947030415532e-15
+ a0 = 1.34374920090936 la0 = -1.50898108050853e-06 wa0 = -2.10741833849894e-07 pa0 = 6.22030879880252e-13
+ keta = 0.0484246926069015 lketa = -2.33742998460202e-07 wketa = -1.74065212117695e-08 pketa = 7.66546407586974e-14
+ a1 = 0.0
+ a2 = 0.5
+ ags = -0.552026352943877 lags = 2.70779171805028e-06 wags = 2.38700357290689e-07 pags = -9.68599281673698e-13
+ b0 = -3.99123276192523e-07 lb0 = 1.19471325457128e-12 wb0 = 1.45226997396837e-13 pb0 = -4.5541696565285e-19
+ b1 = -5.45020871218005e-07 lb1 = 2.36694507299702e-12 wb1 = 2.4931898206934e-13 pb1 = -9.80297146279884e-19
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.135409768368836+0*(0.009/sqrt(l*w*mult))} lvoff = 2.93381891993061e-07 wvoff = -3.66673408725937e-09 pvoff = -1.05121814675205e-13
+ nfactor = {1.36584796581678+0*(0.02/sqrt(l*w*mult))} lnfactor = 2.29770955560247e-06 wnfactor = 6.18948199682681e-09 pnfactor = -9.14475995008673e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.625725e-05 wcit = -3.9446079435e-12
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.61956728893375 leta0 = -2.12239062885735e-06 weta0 = -3.27957524817269e-07 peta0 = 1.29002256365635e-12
+ etab = -1.41587118763606 letab = 5.29399104592239e-06 wetab = 8.05784011556849e-07 petab = -3.16955543837893e-12
+ dsub = 0.728232836085836 ldsub = -6.61744701907814e-07 wdsub = 4.26769677930068e-08 pdsub = -1.67870066198631e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.933071121847248 lpclm = -1.23913990442229e-06 wpclm = -6.81378646670225e-08 ppclm = 1.20262323496339e-12
+ pdiblc1 = 0.283093325998353 lpdiblc1 = 4.20517936718848e-07 wpdiblc1 = -2.80568043827133e-08 ppdiblc1 = 1.10361580323425e-13
+ pdiblc2 = -0.000322105036964595 lpdiblc2 = 6.34122322342542e-09 wpdiblc2 = 5.64891277582616e-10 ppdiblc2 = -2.22200266482761e-15
+ pdiblcb = -0.025
+ drout = 0.549889384665144 ldrout = 3.97701559727329e-08 wdrout = 8.81362128227755e-08 pdrout = -3.46684233819452e-13
+ pscbe1 = 194074124.081267 lpscbe1 = 126.956752564349 wpscbe1 = -12.1436852565825 ppscbe1 = 4.5908692984383e-5
+ pscbe2 = 1.57204815386821e-08 lpscbe2 = -2.88380768374483e-15 wpscbe2 = -1.64947749020831e-16 ppscbe2 = 6.6628465391861e-22
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.67211338883234e-05 lalpha0 = -8.49601506481113e-11 walpha0 = 3.81447746174115e-13 palpha0 = 8.06284082634694e-18
+ alpha1 = -2.176594916125e-10 lalpha1 = 8.56164698555227e-16 walpha1 = 7.62691918179696e-17 palpha1 = -3.00005247361943e-22
+ beta0 = 112.041509626682 lbeta0 = -0.000288917237065567 wbeta0 = -2.5734261884052e-05 pbeta0 = 9.89825342936624e-11
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 6.23647978325198e-08 lagidl = -2.8611333107923e-13 wagidl = -1.19204094422541e-15 pagidl = 1.06785067766999e-19
+ bgidl = 3291941067.20001 lbgidl = -5684.09691775331 wbgidl = -591.970104384086 pbgidl = 0.00196897313911334
+ cgidl = 118.927953447251 lcgidl = 0.00425240230047547 wcgidl = 0.000395074413617083 pcgidl = -1.55402718133486e-9
+ egidl = 1.35687309410667 legidl = -2.2352161603521e-06 wegidl = -5.94817731375635e-08 pegidl = 9.79014143839016e-13
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.4141357500325 lkt1 = -5.97358786568411e-07 wkt1 = -4.57615150907818e-08 pkt1 = 1.80003148417166e-13
+ kt2 = -0.019032
+ at = 1162434.72760696 lat = -2.5413043609734 wat = -0.318280778264086 pat = 8.42984744562323e-7
+ ute = -1.17280632105473 lute = -7.77053209467632e-07 wute = -1.25768285654483e-07 pute = 3.9540691602304e-13
+ ua1 = -4.9057671776e-10 lua1 = 2.01660069867255e-15 wua1 = 1.23259516440783e-32 pua1 = -5.87747175411144e-38
+ ub1 = -7.79729129484788e-19 lub1 = -6.37255686952594e-24 wub1 = -2.95390579910996e-25 pub1 = 1.1619203230328e-30
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.84 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 4.2e-07 wmax = 7.0e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.014/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.7630534664461+0*(0.0/sqrt(l*w*mult))} lvth0 = -2.22463382434544e-07 wvth0 = -1.2304354414697e-07 pvth0 = 1.40877167378904e-13
+ k1 = 0.509824683240378 lk1 = 2.03638085738249e-08 wk1 = 3.1529955777166e-08 pk1 = -1.28374671077905e-14
+ k2 = 0.0644639691695102 lk2 = -1.96822042926467e-08 wk2 = -1.95989352330594e-08 pk2 = 1.40015561632542e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -191819.554779337 lvsat = 0.220560159555659 wvsat = 0.126569581920099 pvsat = -1.03396107051723e-7
+ ua = 1.96280803356906e-09 lua = 4.0090633831424e-16 wua = 2.98591116024205e-17 pua = -1.99430374828155e-22
+ ub = -2.63609312834823e-18 lub = 2.74741542482643e-24 wub = 1.47163625072778e-24 pub = -1.80945150972307e-30
+ uc = 1.65034745632381e-11 luc = -1.62659849297914e-17 wuc = -1.21671371739337e-17 puc = 1.02541744956501e-23
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0087502220290968 lu0 = 8.88660089389433e-09 wu0 = 4.71047259659454e-09 pu0 = -5.827231839404e-15
+ a0 = 0.275198059765772 la0 = 5.57067893648295e-07 wa0 = 2.92597863975298e-07 pa0 = -3.51178942563247e-13
+ keta = -0.0862648743221764 lketa = 2.66799526450044e-08 wketa = 2.82501048000579e-08 pketa = -1.1622673918301e-14
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.881287823868531 lags = -6.35284093873932e-08 wags = -2.82967790514445e-07 pags = 4.0048690448269e-14
+ b0 = -4.06268050822124e-08 lb0 = 5.01558535197134e-13 wb0 = 8.70871748904213e-14 pb0 = -3.43003328137582e-19
+ b1 = 6.17574440477764e-06 lb1 = -1.06276881919669e-11 wb1 = -3.78966418358317e-12 pb1 = 6.82909699942508e-18
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {0.157930960336333+0*(0.009/sqrt(l*w*mult))} lvoff = -2.73793873662026e-07 wvoff = -1.47303867373694e-07 pvoff = 1.72601300719783e-13
+ nfactor = {3.75835699977441+0*(0.02/sqrt(l*w*mult))} lnfactor = -2.32821862409979e-06 wnfactor = -1.12432366499293e-06 pnfactor = 1.27137682726176e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.625725e-05 wcit = -3.9446079435e-12
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -0.66455268476794 leta0 = 3.60461760894735e-07 weta0 = 4.70820729392552e-07 peta0 = -2.54419184749606e-13
+ etab = 2.56461756258936 letab = -2.40230385508222e-06 wetab = -1.61419585297655e-06 petab = 1.50948772959573e-12
+ dsub = 0.395694935345119 ldsub = -1.87810081361348e-08 wdsub = -5.02680860929151e-08 pdsub = 1.18396602150683e-14
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.759193736086849 lpclm = 2.03286265971758e-06 wpclm = 1.21665428887037e-06 ppclm = -1.28152881786192e-12
+ pdiblc1 = 0.310368282569688 lpdiblc1 = 3.67781671813389e-07 wpdiblc1 = 1.48934386705293e-07 ppdiblc1 = -2.31851772601192e-13
+ pdiblc2 = 0.00282037628669519 lpdiblc2 = 2.65219871722617e-10 wpdiblc2 = -4.97845289622765e-10 ppdiblc2 = -1.67196198453168e-16
+ pdiblcb = -0.025
+ drout = 1.23125700855358 ldrout = -1.27765755165368e-06 wdrout = -5.07738750173048e-07 pdrout = 8.05442986507788e-13
+ pscbe1 = 278590340.728144 lpscbe1 = -36.4557749034709 wpscbe1 = -0.286072397766247 ppscbe1 = 2.29819392337974e-5
+ pscbe2 = 1.43949464126998e-08 lpscbe2 = -3.20878889982371e-16 wpscbe2 = 7.50312923575879e-17 ppscbe2 = 2.02283977518229e-22
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -1.65365575573375e-06 lalpha0 = -1.07623029973787e-11 walpha0 = 1.04253755094909e-12 palpha0 = 6.78462038336551e-18
+ alpha1 = 2.25145e-10 walpha1 = -7.889215887e-17
+ beta0 = -31.6142536658918 lbeta0 = -1.11581004605592e-05 wbeta0 = 2.18210331965002e-05 pbeta0 = 7.03413347893928e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -1.0734088475985e-07 lagidl = 4.20134547415294e-14 wagidl = 6.7734908671518e-14 pagidl = -2.64855339497886e-20
+ bgidl = 604399922.244534 lbgidl = -487.722676276179 wbgidl = 267.355233617512 pbgidl = 0.000307463301460561
+ cgidl = 3561.32942770907 lcgidl = -0.00240349816201712 wcgidl = -0.000794523412985263 pcgidl = 7.46066164389905e-10
+ egidl = -0.631385398678168 legidl = 1.60909157673986e-06 wegidl = 9.7149312910747e-07 pegidl = -1.01438098452627e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.783835211277 lkt1 = 1.17456970245136e-07 wkt1 = 8.56313322002886e-08 pkt1 = -7.40455787843552e-14
+ kt2 = -0.019032
+ at = -345100.8496167 lat = 0.373523215266438 wat = 0.242316513338009 pat = -2.40932921736786e-7
+ ute = -1.69128454625855 lute = 2.25427031355088e-07 wute = 1.52233306868667e-07 pute = -1.42110553128435e-13
+ ua1 = 5.524e-10
+ ub1 = -3.71612072711668e-18 lub1 = -6.95029033546699e-25 wub1 = 7.89398976987143e-26 pub1 = 4.3815047292204e-31
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.81e-6
+ sbref = 2.81e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.85 pmos
* DC IV MOS Parameters
+ lmin = 8.0e-07 lmax = 1e-06 wmin = 4.2e-07 wmax = 7.0e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.02/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.45586106088675+0*(0.0/sqrt(l*w*mult))} lvth0 = 4.24275971013772e-07 wvth0 = 3.08026268729442e-07 pvth0 = -2.61528658290292e-13
+ k1 = 0.271348711926804 lk1 = 2.42982320174903e-07 wk1 = 1.81866638949071e-07 pk1 = -1.5317751253218e-13
+ k2 = 0.0708341635851132 lk2 = -2.56288126305841e-08 wk2 = -2.71818738776096e-08 pk2 = 2.1080267302635e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -75927.1805401669 lvsat = 0.112374048741523 wvsat = 0.0711832592642172 pvsat = -5.16926979208441e-8
+ ua = 1.57443646651291e-09 lua = 7.63453138018992e-16 wua = 3.50962497163485e-16 pua = -4.99181990766338e-22
+ ub = 4.19880401539501e-18 lub = -3.63299523334362e-24 wub = -3.28774201688561e-24 pub = 2.63345189998537e-30
+ uc = -1.19401376134007e-12 luc = 2.5470890864395e-19 wuc = -1.01053434918965e-18 puc = -1.60570024262597e-25
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0293506461972199 lu0 = -1.03439980691694e-08 wu0 = -8.45598667842814e-09 pu0 = 6.46372372612606e-15
+ a0 = 1.47735418590846 la0 = -5.65150860886531e-07 wa0 = -4.65248570881806e-07 pa0 = 3.56274493608034e-13
+ keta = -0.135851375848699 lketa = 7.29691997525206e-08 wketa = 6.50764179112747e-08 pketa = -4.60002213391875e-14
+ a1 = 0.0
+ a2 = 0.5
+ ags = 2.08839431425812 lags = -1.19036835369853e-06 wags = -1.04393496469499e-06 pags = 7.50415352381675e-13
+ b0 = 2.31816604759431e-06 lb0 = -1.70038638674067e-12 wb0 = -1.30853507470749e-12 pb0 = 9.59817019973321e-19
+ b1 = -2.43129995569249e-05 lb1 = 1.78337067400022e-11 wb1 = 1.64571326786463e-11 pb1 = -1.20713891054505e-17
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.511681296868581+0*(0.009/sqrt(l*w*mult))} lvoff = 3.51292516500047e-07 wvoff = 2.74823717241826e-07 pvoff = -2.21456910156729e-13
+ nfactor = {-1.00748760227795+0*(0.02/sqrt(l*w*mult))} lnfactor = 2.1207211411391e-06 wnfactor = 1.71131065163115e-06 pnfactor = -1.3757019854784e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.625725e-05 wcit = -3.9446079435e-12
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.651279849052799 leta0 = -8.67874488589594e-07 weta0 = -3.87806133455979e-07 peta0 = 5.47113284853812e-13
+ etab = -0.00528913092795897 letab = -3.28310715033347e-09 wetab = 5.978965475709e-10 petab = 2.06969044621312e-15
+ dsub = 1.29757492496141 ldsub = -8.60690487842888e-07 wdsub = -6.1881864282696e-07 pdsub = 5.42584447679083e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.51924218586239 lpclm = -9.40686656016465e-08 wpclm = -2.19685386941967e-07 ppclm = 5.93014512072721e-14
+ pdiblc1 = 0.61751200219404 lpdiblc1 = 8.10614738254593e-08 wpdiblc1 = -4.46908570082157e-08 ppdiblc1 = -5.11016394684126e-14
+ pdiblc2 = 0.0275178249026702 lpdiblc2 = -2.27899718985331e-08 wpdiblc2 = -1.60672650818251e-08 ppdiblc2 = 1.43669350246667e-14
+ pdiblcb = -0.025
+ drout = -1.81310380165778 ldrout = 1.56426848648268e-06 wdrout = 1.41144457074906e-06 pdrout = -9.86124239489601e-13
+ pscbe1 = 239227545.331441 lpscbe1 = 0.289591413328253 wpscbe1 = 24.5284699970875 ppscbe1 = -1.82560164510635e-7
+ pscbe2 = 1.20179400727454e-08 lpscbe2 = 1.89806841339669e-15 wpscbe2 = 1.57351035110284e-15 ppscbe2 = -1.19655371621576e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -6.15303613206746e-05 lalpha0 = 4.51329010310214e-11 walpha0 = 3.87891719993212e-11 palpha0 = -2.84520516073621e-17
+ alpha1 = 6.84117416125e-10 lalpha1 = -4.28453045314768e-16 walpha1 = -3.68231123829697e-16 palpha1 = 2.70099370484702e-22
+ beta0 = -214.353396644688 lbeta0 = 0.000159429803205862 wbeta0 = 0.000137020885365191 pbeta0 = -1.00505504519794e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 2.83909703840722e-06 lagidl = -2.70850107872455e-12 wagidl = -1.79002797352098e-12 pagidl = 1.70774540539132e-18
+ bgidl = -790894130.616993 lbgidl = 814.791298540321 wbgidl = 1146.95697630574 pbgidl = -0.000513649323347609
+ cgidl = 22779.5546494472 lcgidl = -0.0203438074976358 wcgidl = -0.0137337065399794 pcgidl = 1.28248583093546e-8
+ egidl = 6.76649370428809 legidl = -5.29686555527466e-06 wegidl = -3.69217424467708e-06 pegidl = 3.33917582723848e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.5588714309525 lkt1 = -9.25478435066862e-08 wkt1 = -5.7343199581533e-08 pkt1 = 5.94218615066339e-14
+ kt2 = -0.019032
+ at = 220173.983225 lat = -0.154163667565454 wat = -0.0736462247659393 pat = 5.40198740969403e-8
+ ute = -1.33977425 lute = -1.02709587753751e-7
+ ua1 = 5.524e-10
+ ub1 = -4.46065775e-18 wub1 = 5.48300504146502e-25
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.41e-6
+ sbref = 2.41e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.86 pmos
* DC IV MOS Parameters
+ lmin = 6e-07 lmax = 8.0e-07 wmin = 4.2e-07 wmax = 7.0e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.02/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.594966578964661+0*(0.0/sqrt(l*w*mult))} lvth0 = -2.07194435948487e-07 wvth0 = -1.47295168605556e-07 pvth0 = 7.24518926021155e-14
+ k1 = 0.566868317130449 lk1 = 2.62172121600024e-08 wk1 = -2.2676311140816e-08 pk1 = -3.14423592649724e-15
+ k2 = 0.0390698858818645 lk2 = -2.32955611386267e-09 wk2 = 3.80135079961148e-09 pk2 = -1.64608291423005e-15
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 165284.918813144 lvsat = -0.0645562321946272 wvsat = -0.0350647532106668 pvsat = 2.62407504695457e-8
+ ua = 1.13538349967831e-08 lua = -6.40978458092681e-15 wua = -2.91980146646404e-15 pua = 1.89993973037427e-21
+ ub = -1.36955562966192e-17 lub = 9.49260752732037e-24 wub = 4.31974738187873e-24 pub = -2.94667961145527e-30
+ uc = -1.57743823857139e-12 luc = 5.35952679815508e-19 wuc = -6.8793565957958e-19 puc = -3.97197776085032e-25
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0218502812921967 lu0 = -4.8424429095104e-09 wu0 = -6.58863636163366e-10 pu0 = 7.44494989009622e-16
+ a0 = -0.159492774280233 la0 = 6.35484568646673e-07 wa0 = 4.4728473529021e-07 pa0 = -3.1307324913567e-13
+ keta = 0.242438022065408 lketa = -2.04507965064466e-07 wketa = -1.05226460830984e-07 pketa = 7.89177917326533e-14
+ a1 = 0.0
+ a2 = 0.5
+ ags = -2.57748979023929 lags = 2.23208096637085e-06 wags = 1.02067710557998e-06 pags = -7.63987924225361e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {0.152511819939713+0*(0.009/sqrt(l*w*mult))} lvoff = -1.35896455644421e-07 wvoff = -9.08097913919269e-08 pvoff = 4.67370965936727e-14
+ nfactor = {3.99103946874982+0*(0.02/sqrt(l*w*mult))} lnfactor = -1.54572345809512e-06 wnfactor = -8.62314331499984e-07 pnfactor = 5.120648077732e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 6.29776166125e-05 lcit = -3.42696225121018e-11 wcit = -2.49892885524697e-11 pcit = 1.54363784500823e-17
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -1.76089012645047 leta0 = 9.01464249291929e-07 weta0 = 1.15844805881684e-06 peta0 = -5.87071896449261e-13
+ etab = -0.155644488644474 letab = 1.07003299511519e-07 wetab = 8.80833919068215e-08 petab = -6.2101357827274e-14
+ dsub = -0.307176865581564 ldsub = 3.16402974279334e-07 wdsub = 4.35615195718986e-07 pdsub = -2.30848045063561e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.44967663601925 lpclm = -4.30419869639547e-08 wpclm = -2.57523793113786e-07 ppclm = 8.70561113263325e-14
+ pdiblc1 = 0.251566651892491 lpdiblc1 = 3.49484217998397e-07 wpdiblc1 = 9.70297007678191e-08 ppdiblc1 = -1.55054377199923e-13
+ pdiblc2 = -0.0295108219662219 lpdiblc2 = 1.90408257230335e-08 wpdiblc2 = 1.56549998984857e-08 ppdiblc2 = -8.90150494971618e-15
+ pdiblcb = -0.025
+ drout = -2.43206044796381 ldrout = 2.01827628133138e-06 wdrout = 8.37587562449697e-07 pdrout = -5.6519725461698e-13
+ pscbe1 = -238232807.248289 lpscbe1 = 350.509147332324 wpscbe1 = 120.593867402296 ppscbe1 = -7.06470094882183e-5
+ pscbe2 = 1.26874550366343e-08 lpscbe2 = 1.40697583980944e-15 wpscbe2 = 1.20882110364447e-15 ppscbe2 = -9.29052329758809e-22
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -0.000139543517050514 lalpha0 = 1.02355940824637e-10 walpha0 = 3.03441987019897e-11 palpha0 = -2.2257621468903e-17
+ alpha1 = 3.667525e-10 lalpha1 = -1.956642925125e-16
+ beta0 = -135.762188071794 lbeta0 = 0.000101782758761602 wbeta0 = 9.28162801003437e-06 pbeta0 = -6.80812055350026e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -3.03775285053067e-06 lagidl = 1.60219769906084e-12 wagidl = 1.86663725906941e-12 pagidl = -9.74436826039896e-19
+ bgidl = -4003043496.14053 lbgidl = 3170.91891889866 wbgidl = 1974.26276368814 pbgidl = -0.00112048225492154
+ cgidl = -16608.9958969678 lcgidl = 0.00854789127091236 wcgidl = 0.0114234079636489 pcgidl = -5.62801096462931e-9
+ egidl = -2.92307863127995 legidl = 1.81048420072618e-06 wegidl = 2.34288649702247e-06 pegidl = -1.08757140210185e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.9026161753375 lkt1 = 1.59590645223433e-07 wkt1 = 8.68016894879086e-08 pkt1 = -4.63091353502468e-14
+ kt2 = -0.019032
+ at = 10000.0
+ ute = -1.515691548875 lute = 2.63266305575581e-08 wute = -2.10446806089696e-07 pute = 1.54363784500823e-13
+ ua1 = 5.5346701e-10 lua1 = -7.82657170049756e-19
+ ub1 = -1.13723690745687e-17 lub1 = 5.0697748151278e-24 wub1 = 2.01090580646989e-24 pub1 = -1.07282830228072e-30
+ uc1 = -5.4204995714961e-10 luc1 = 3.17497607819025e-16 wuc1 = 1.51673222084966e-16 puc1 = -1.11253066765433e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.02e-6
+ sbref = 2.01e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.87 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 6e-07 wmin = 4.2e-07 wmax = 7.0e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.32475e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 3.4797e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.22435e-08+0*(1.22435e-08*(0.02/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.858939541650637+0*(0.0/sqrt(l*w*mult))} lvth0 = -6.63635404907059e-08 wvth0 = -1.00881151410344e-07 pvth0 = 4.76897823583839e-14
+ k1 = 0.828121187608434 lk1 = -1.13162500504354e-07 wk1 = -5.72084084154473e-08 pk1 = 1.52788106300048e-14
+ k2 = -0.0517585496340073 lk2 = 4.61278683760325e-08 wk2 = 1.38412360274919e-08 pk2 = -7.00241188273043e-15
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -49491.0128020305 lvsat = 0.0500278012017265 wvsat = 0.0365401530218655 pvsat = -1.19608250300415e-8
+ ua = -8.58728448262606e-09 lua = 4.22890236693535e-15 wua = 1.33299563854766e-15 pua = -3.68948789134998e-22
+ ub = 9.23324872200117e-18 lub = -2.7400245941387e-24 wub = 7.58908664463572e-25 pub = -1.04695435152069e-30
+ uc = 8.38330237750654e-12 luc = -4.77815224256515e-18 wuc = -9.46786450052378e-19 puc = -2.59099585113845e-25
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = -0.00822659735566295 lu0 = 1.1203722233516e-08 wu0 = 8.1939535678444e-09 pu0 = -3.97852725341454e-15
+ a0 = -1.02942320271472 la0 = 1.09959680186861e-06 wa0 = 1.50928195270064e-06 pa0 = -8.79654074610223e-13
+ keta = -0.332281138624689 lketa = 1.02107580759504e-07 wketa = 9.40672612276702e-08 pketa = -2.74064054542492e-14
+ a1 = 0.0
+ a2 = 0.5
+ ags = -0.951222773410365 lags = 1.36445938155753e-06 wags = 1.10520651179226e-06 pags = -8.09084785086648e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0186024814734855+0*(0.009/sqrt(l*w*mult))} lvoff = -4.46061202689723e-08 wvoff = -7.78533519393647e-08 pvoff = 3.98247713635335e-14
+ nfactor = {1.28139824631473+0*(0.02/sqrt(l*w*mult))} lnfactor = -1.00116317719892e-07 wnfactor = -6.57199099627246e-07 pnfactor = 4.02634805992935e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -5.00579916125e-05 lcit = 2.60354396539768e-11 wcit = 2.10446806089697e-11 pcit = -9.12297426739141e-18
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -1.02223390386524 leta0 = 5.07387461261599e-07 weta0 = 5.28285490733458e-07 peta0 = -2.50877015563937e-13
+ etab = 0.166548288985837 letab = -6.48881583181401e-08 wetab = -9.30442376434748e-08 petab = 3.45311381759568e-14
+ dsub = 0.411800130378045 ldsub = -6.71748479500968e-08 wdsub = -1.95067496792489e-08 pdsub = 1.19617884161241e-14
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 3.08622371844746 lpclm = -9.16148038174815e-07 wpclm = -6.84601969442357e-07 ppclm = 3.14904453788507e-13
+ pdiblc1 = 5.18359751374971 lpdiblc1 = -2.28177890695674e-06 wpdiblc1 = -1.74453450561682e-06 ppdiblc1 = 8.27429334727312e-13
+ pdiblc2 = 0.0346610542328155 lpdiblc2 = -1.51951910885339e-08 wpdiblc2 = -1.66887748925185e-08 ppdiblc2 = 8.35406062015852e-15
+ pdiblcb = -0.025
+ drout = 1.93165661226968 ldrout = -3.09788588888486e-07 wdrout = -5.90256990801699e-07 pdrout = 1.96564953765407e-13
+ pscbe1 = 295567458.616102 lpscbe1 = 65.7240364923409 wpscbe1 = 65.8349006836572 ppscbe1 = -4.14328269489906e-5
+ pscbe2 = 1.76299178337874e-08 lpscbe2 = -1.22985277478578e-15 wpscbe2 = -2.70063105039295e-15 ppscbe2 = 1.15665994168093e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.000148951944115215 lalpha0 = -5.15578301845848e-11 walpha0 = -3.17667230235045e-11 palpha0 = 1.08788658262568e-17
+ alpha1 = 0.0
+ beta0 = 74.1016569160298 lbeta0 = -1.01806518586276e-05 wbeta0 = -7.64359079777457e-06 pbeta0 = 2.22156830655985e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -2.8380720443785e-07 lagidl = 1.3295392714209e-13 wagidl = 1.86053928846617e-13 pagidl = -7.78372164493835e-20
+ bgidl = 2004034644.7951 lbgidl = -33.8873046812005 wbgidl = -284.886346654748 pbgidl = 8.47850911919433e-5
+ cgidl = -7163.23118513063 lcgidl = 0.00350852856832367 wcgidl = 0.00491075505728146 pcgidl = -2.15347807581774e-9
+ egidl = -0.306521566937207 legidl = 4.14537924114001e-07 wegidl = 8.59743979336721e-07 pegidl = -2.96307453203915e-13
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.413827848322501 lkt1 = -1.01180371180705e-07 wkt1 = 3.42001453309396e-09 pkt1 = -1.82459485347824e-15
+ kt2 = -0.019032
+ at = 102201.5281925 lat = -0.0491899762983397 wat = -0.0444601889302212 pat = 2.37197330952177e-8
+ ute = -1.846678704328 lute = 2.0290993292751e-07 wute = 3.96269507541117e-07 pute = -1.69322402402784e-13
+ ua1 = 5.52e-10
+ ub1 = 4.66937241668996e-19 lub1 = -1.24655430111662e-24 wub1 = 7.37355133335053e-25 pub1 = -3.93382650409918e-31
+ uc1 = 1.12380077112576e-09 luc1 = -5.71242084969527e-16 wuc1 = -5.34895108118525e-16 puc1 = 2.5503457023978e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 2.36876351e-10
+ cgso = 2.36876351e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 1.19869905e-11
+ cgdl = 1.19869905e-11
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 3.28555e-8
+ dwc = 2.252e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.000818818773
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 1.040674614e-10
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.539132e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 1.81e-6
+ sbref = 1.81e-6
+ wlod = {0+0.0}
+ kvth0 = {0+3.5e-8}
+ lkvth0 = {0+0.0}
+ wkvth0 = {0+6.5e-7}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+7.0e-8}
+ lku0 = {0+0.0}
+ wku0 = {0+0.0}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+0.4}
+ steta0 = 0.0
+ tku0 = 0.0
.ends sky130_fd_pr__pfet_g5v0d10v5
