** NGSPICE Simulation bench



.GLOBAL
** Default values that can be modified in the corners
.PARAM vdd=3.3 vcm=1.65 c1=6p ib=100u
.TEMP 25.0
**
** Process, Voltage and Temperature settings for nominal.
** Pyhton script replaces this include to simulate other corners
**
.lib "../device_models/ptm130/ptm-130.lib" FF
**
** Design variables for the circuit being simulated
**
.include 'design_var.inc'

*********** Unit Under Test ********************
.include "ssvcamp.cir"

*********** Test-bench *************************
mnmbias halfvdd halfvdd 0 0 nmos33 w='_w10/_nf10' l='_l10'  m='_nf10'
g2 cmfb 0 VCCS halfvdd 0 -1
g1 cmfb 0 VCCS outputn 0 -500m
g0 cmfb 0 VCCS outputp 0 -500m
e3 output 0 VCVS outputp outputn 1
i0 cmfb 0 DC 'vcm'
xinova cmfb 0 vddnet in_n in_p outputn outputp ssvcamp
cload2 outputp 0 'c1'
cload1 outputn 0 'c1'
r0 cmfb 0 1
cload3 output 0 'c1'
ibias vddnet halfvdd DC 'ib'
vin in_n 0 DC 'vcm'
vip in_p 0 DC 'vcm' AC 1 sin 'vcm' 100e-3 1e3
vdc vddnet 0 DC 'vdd'
************************************************

*********** OPTIONS ****************************
.OPTION KEEPOPINFO
************************************************


************************************************
** make params acessible in control
.csparam ib = {ib}
.csparam c1 = {c1}
************************************************
.control
set units = degrees

***********************************************
** Run OP and save dc current, deltas and
** overdrives.

OP 
let idd = mag(i(vdc))  
print idd
** Overdrive and delta for  PMOS
let   vov_mpm0 = @m.xinova.mpm0[vth]   - @m.xinova.mpm0[vgs] 
let delta_mpm0 = @m.xinova.mpm0[vdsat] - @m.xinova.mpm0[vds]
print vov_mpm0 delta_mpm0 

let   vov_mpm1 = @m.xinova.mpm1[vth]   - @m.xinova.mpm1[vgs] 
let delta_mpm1 = @m.xinova.mpm1[vdsat] - @m.xinova.mpm1[vds]
print vov_mpm1 delta_mpm1 

let   vov_mpm2 = @m.xinova.mpm2[vth]   - @m.xinova.mpm2[vgs] 
let delta_mpm2 = @m.xinova.mpm2[vdsat] - @m.xinova.mpm2[vds]
print vov_mpm2 delta_mpm2 

let   vov_mpm3 = @m.xinova.mpm3[vth]   - @m.xinova.mpm3[vgs] 
let delta_mpm3 = @m.xinova.mpm3[vdsat] - @m.xinova.mpm3[vds]
print vov_mpm3 delta_mpm3 

** Overdrive and delta for NMOS
let   vov_mnm4 = @m.xinova.mnm4[vgs] - @m.xinova.mnm4[vth] 
let delta_mnm4 = @m.xinova.mnm4[vds] - @m.xinova.mnm4[vdsat]
print vov_mnm4 delta_mnm4

let   vov_mnm5 = @m.xinova.mnm5[vgs] - @m.xinova.mnm5[vth] 
let delta_mnm5 = @m.xinova.mnm5[vds] - @m.xinova.mnm5[vdsat]
print vov_mnm5 delta_mnm5

let   vov_mnm6 = @m.xinova.mnm6[vgs] - @m.xinova.mnm6[vth] 
let delta_mnm6 = @m.xinova.mnm6[vds] - @m.xinova.mnm6[vdsat]
print vov_mnm6 delta_mnm6

let   vov_mnm7 = @m.xinova.mnm7[vgs] - @m.xinova.mnm7[vth] 
let delta_mnm7 = @m.xinova.mnm7[vds] - @m.xinova.mnm7[vdsat]
print vov_mnm7 delta_mnm7

let   vov_mnm8 = @m.xinova.mnm8[vgs] - @m.xinova.mnm8[vth] 
let delta_mnm8 = @m.xinova.mnm8[vds] - @m.xinova.mnm8[vdsat]
print vov_mnm8 delta_mnm8

let   vov_mnm9 = @m.xinova.mnm9[vgs] - @m.xinova.mnm9[vth] 
let delta_mnm9 = @m.xinova.mnm9[vds] - @m.xinova.mnm9[vdsat]
print vov_mnm9 delta_mnm9

let   vov_mnm10 = @m.xinova.mnm10[vgs] - @m.xinova.mnm10[vth] 
let delta_mnm10 = @m.xinova.mnm10[vds] - @m.xinova.mnm10[vdsat]
print vov_mnm10 delta_mnm10

let   vov_mnm11 = @m.xinova.mnm7[vgs] - @m.xinova.mnm7[vth] 
let delta_mnm11 = @m.xinova.mnm7[vds] - @m.xinova.mnm7[vdsat]
print vov_mnm11 delta_mnm11
************************************************

************************************************
* Run AC
AC DEC 20 1 10G

let vdb_out = vdb(output)
let vp_out = vp(output)

print frequency vdb_out vp_out


************************************************
* Run noise
NOISE V(output, 0) vip dec 20 0.01 10G
print inoise_total onoise_total
print noise2.all

quit

.endc

.END
